--------------------------------------------------------------------------------
--
--
--          **  **     **  ******  ********  ********  ********  **    **
--         **    **   **  **   ** ********  ********  ********  **    **
--        **     *****   **   **    **     **        **        **    **
--       **       **    ******     **     ****      **        ********
--      **       **    **  **     **     **        **        **    **
--     *******  **    **   **    **     ********  ********  **    **
--    *******  **    **    **   **     ********  ********  **    **
--
--                       L Y R T E C H   R D   I N C
--
--------------------------------------------------------------------------------
-- File        : $Id: dsp_mult16x16_16_p.vhd,v 1.1 2010/07/29 14:27:02 francois.blackburn Exp $
--------------------------------------------------------------------------------
-- Description : ADAC250Wrapper
--
--
--------------------------------------------------------------------------------
-- Notes / Assumptions :
--
--------------------------------------------------------------------------------
-- Copyright (c) 2009 Lyrtech RD inc.
-- TODO = legal notice
--------------------------------------------------------------------------------
-- $Log: dsp_mult16x16_16_p.vhd,v $
-- Revision 1.1  2010/07/29 14:27:02  francois.blackburn
-- first commit
--
-- Revision 1.2  2010/07/26 18:08:48  patrick.gilbert
-- work with 31 bit data port
--
-- Revision 1.1  2010/06/17 15:40:21  francois.blackburn
-- first commit
--

--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

package dsp_mult16x16_16_p is

  component dsp_mult16x16_16 IS
    port (
    clk: in std_logic;
    a: in std_logic_vector(15 downto 0);
    b: in std_logic_vector(15 downto 0);
    p: out std_logic_vector(31 downto 0));
  end component;

end dsp_mult16x16_16_p;

