--------------------------------------------------------------------------------
--
--    ****                              *
--   ******                            ***
--   *******                           ****
--   ********    ****  ****     **** *********    ******* ****    ***********
--   *********   ****  ****     **** *********  **************  *************
--   **** *****  ****  ****     ****   ****    *****    ****** *****     ****
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      ****
--  ****    *********  ****     ****   ****   ****       ****  ****      ****
--  ****     ********  ****    *****  ****    *****     *****  ****      ****
--  ****      ******   ***** ******   *****    ****** *******  ****** *******
--  ****        ****   ************    ******   *************   *************
--  ****         ***     ****  ****     ****      *****  ****     *****  ****
--                                                                       ****
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       ****
--                                                                        ***
--
--------------------------------------------------------------------------------
-- File        : $Id: Bustestin_wrapper_p.vhd,v 1.1 2013/02/07 14:46:12 julien.roy Exp $
--------------------------------------------------------------------------------
-- Description : Bustestin_wrapper_p
--
--
--------------------------------------------------------------------------------
-- Notes / Assumptions :
--
--------------------------------------------------------------------------------
-- Copyright (c) 2013 Nutaq inc.
--------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

Package Bustestin_wrapper_p is

  component Bustestin_wrapper is
    PORT (
      clk           : IN  std_logic;
      ce            : IN  std_logic;
      start         : IN  std_logic;
      nRstErr       : IN  std_logic;
      pattern       : IN std_logic_vector(13 DOWNTO 0);
      lock          : OUT std_logic;
      errorCnt      : OUT std_logic_vector(31 DOWNTO 0);
      dataCountDiv1024 : out std_logic_vector(31 downto 0);
      errorMask     : OUT std_logic_vector(13 DOWNTO 0)
    );
  end component;

end Bustestin_wrapper_p;