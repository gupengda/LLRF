--------------------------------------------------------------------------------
--
--
--          **  **     **  ******  ********  ********  ********  **    **
--         **    **   **  **   ** ********  ********  ********  **    **
--        **     *****   **   **    **     **        **        **    **
--       **       **    ******     **     ****      **        ********
--      **       **    **  **     **     **        **        **    **
--     *******  **    **   **    **     ********  ********  **    **
--    *******  **    **    **   **     ********  ********  **    **
--
--                       L Y R T E C H   R D   I N C
--
--------------------------------------------------------------------------------
-- File        : $Id: lyt_mestor_mbb1_e.vhd,v 1.4 2011/02/21 22:00:23 francois.blackburn Exp $
--------------------------------------------------------------------------------
-- Description : I/O ring file.
--               Generated by generate_ioring_v2.pl (2.06)
--
--------------------------------------------------------------------------------
-- Notes / Assumptions :
--
--------------------------------------------------------------------------------
-- Copyright (c) 2010 Lyrtech RD inc.
--------------------------------------------------------------------------------
-- $Log: lyt_mestor_mbb1_e.vhd,v $
-- Revision 1.4  2011/02/21 22:00:23  francois.blackburn
-- change core name
--
-- Revision 1.3  2010/09/29 21:27:34  francois.blackburn
-- fix bit shift bug
--
-- Revision 1.2  2010/06/18 14:19:43  francois.blackburn
-- change LYR for lyt
--
-- Revision 1.1  2010/04/01 17:55:15  francois.blackburn
-- first commit
--
--------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;

library UNISIM;
  use UNISIM.vcomponents.all;

entity lyt_mestor_mbb1 is
port
(
    -- User Ports
    i_SysClk_p                 : in std_logic;
    i_Reset_p                  : in std_logic;
    o_DelayRdy_p               : out std_logic;
    iv32_GpioDIn_p             : in std_logic_vector(31 downto 0);
    iv32_GpioDir_p             : in std_logic_vector(31 downto 0);
    ov32_GpioDOut_p            : out std_logic_vector(31 downto 0);
    i_SetGpioDir_p             : in std_logic;
    o_SetGpioDirAck_p          : out std_logic;
    i_Start_p                  : in std_logic;
    o_StartAck_p               : out std_logic;
    ov12_AdcData0_p            : out std_logic_vector(11 downto 0);
    ov12_AdcData1_p            : out std_logic_vector(11 downto 0);
    ov12_AdcData2_p            : out std_logic_vector(11 downto 0);
    ov12_AdcData3_p            : out std_logic_vector(11 downto 0);
    o_AdcData0Valid_p          : out std_logic;
    o_AdcData1Valid_p          : out std_logic;
    o_AdcData2Valid_p          : out std_logic;
    o_AdcData3Valid_p          : out std_logic;
    
    
    -- Perseus to Mestor Ports
    odp_DpioSetDir_p           : out std_logic;
    odn_DpioSetDir_p           : out std_logic;
    odp_DpioReset_p            : out std_logic;
    odn_DpioReset_p            : out std_logic;
    odp_DpioConfig_p           : out std_logic;
    odn_DpioConfig_p           : out std_logic;
    idp_DpioResetAck_p         : in std_logic;
    idn_DpioResetAck_p         : in std_logic;
    ov4dp_Dpio_p               : out std_logic_vector(3 downto 0);
    ov4dn_Dpio_p               : out std_logic_vector(3 downto 0);
    iv4dp_Dpio_p               : in std_logic_vector(3 downto 0);
    iv4dn_Dpio_p               : in std_logic_vector(3 downto 0);
    odp_DpioClk_p              : out std_logic;
    odn_DpioClk_p              : out std_logic;
    iv2dp_AdcData_p            : in std_logic_vector(1 downto 0);
    iv2dn_AdcData_p            : in std_logic_vector(1 downto 0)
  );

end entity lyt_mestor_mbb1;
