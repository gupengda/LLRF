--------------------------------------------------------------------------------
--
--    ****                              *
--   ******                            ***
--   *******                           ****
--   ********    ****  ****     **** *********    ******* ****    ***********
--   *********   ****  ****     **** *********  **************  *************
--   **** *****  ****  ****     ****   ****    *****    ****** *****     ****
--   ****  ***** ****  ****     ****   ****   *****      ****  ****      ****
--  ****    *********  ****     ****   ****   ****       ****  ****      ****
--  ****     ********  ****    *****  ****    *****     *****  ****      ****
--  ****      ******   ***** ******   *****    ****** *******  ****** *******
--  ****        ****   ************    ******   *************   *************
--  ****         ***     ****  ****     ****      *****  ****     *****  ****
--                                                                       ****
--          I N N O V A T I O N  T O D A Y  F O R  T O M M O R O W       ****
--                                                                        ***
--
--------------------------------------------------------------------------------
-- Filename:          user_logic.vhd
-- Version:           v1_00_a
-- Description:       User Logic implementation module
-- Generated by:      khalid.bensadek
-- Date:              2012-09-21 10:41:46
-- Generated:         using Nutaq REGGENUTIL based on Xilinx IPIF Wizard.
-- VHDL Standard:     VHDL'93
--------------------------------------------------------------------------------
-- Copyright (c) 2012 Nutaq inc.
--------------------------------------------------------------------------------
-- Register Memory Map & Description
--------------------------------------------------------------------------------
-- BASEADDR + 0x0   COREID    Core ID
--   31:0 coreId R

-- BASEADDR + 0x4   BOARDCONTROL    Tx control signal
--   0:0 TxEnable R W O=o_TxEnable_p
--   1:1 RxEnable R W O=o_RxEnable_p
--   11:10 ClkMuxSout R W O=ov2_ClkMuxSout_p
--   12:12 ClkMuxLoad R W O=o_ClkMuxLoad_p
--   13:13 ClkMuxConfig R W O=o_ClkMuxConfig_p
--   14:14 PLLLock R I=i_PLLLock_p
--   15:15 ovrAdcI R I=i_ovrAdcI_p
--   16:16 ovrAdcQ R I=i_ovrAdcQ_p
--   17:17 ovrDacI R I=i_ovrDacI_p
--   18:18 ovrDacQ R I=i_ovrDacQ_p
--   19:19 fmcPps R I=i_fmcPps_p
--   2:2 LimeReset R W O=o_LimeReset_p
--   20:20 ResetOvr R W O=o_ResetOvr_p
--   24:21 rsvd2 R
--   25:25 DesignClkEn R W O=o_DesignClkEn_p
--   26:26 CoreResetPulse P O=o_CoreResetPulse_p
--   27:27 RstFifo R W O=o_RstFifo_p
--   31:28 rsvd3 R
--   7:3 FpgaControl R W O=ov5_FpgaControl_p
--   9:8 ClkMuxSin R W O=ov2_ClkMuxSin_p

-- BASEADDR + 0x8   DACDATAOUTCTRL    DAC data source ctrl
--   23:0 ddsfreq R W O=ov24_ddsfreq_p
--   26:24 dacOutSel R W O=ov3_dacOutSel_p
--   31:27 rsvd0 R

-- BASEADDR + 0xc   LIMESPIDATA    Spi Register to control Lime SPI
--   15:0 limeSpiDataIn W O=ov16_limeSpiDataIn_p  / R iv16_limeSpiDataOut_p
--   31:16 rsvd R

-- BASEADDR + 0x10   TXGAINSPIDATA    Spi Register to control TX gain
--   31:6 rsvd R
--   5:0 txGainSpiData R W O=ov6_txGainSpiData_p

-- BASEADDR + 0x14   RXGAINSPIDATA    Spi Register to control RX gain
--   31:6 rsvd R
--   5:0 rxGainSpiData R W O=ov6_rxGainSpiData_p

-- BASEADDR + 0x18   PLLCTRLSPIDATA    Spi Register to control PLL and GPIO
--   31:0 pllCtrlSpiDataIn R W O=ov32_pllCtrlSpiDataIn_p

-- BASEADDR + 0x1c   REFDACSPIDATA    Spi Register to control reference DAC
--   15:0 refDacSpiData W O=ov16_refDacSpiData_p / R iv16_refDacSpiData_p
--   31:16 rsvd R

-- BASEADDR + 0x20   SPICTRL    control flag of SPI reg.
--   0:0 limeSpiStart R W O=o_limeSpiStart_p
--   1:1 limeSpiBusy R I=i_limeSpiBusy_p
--   10:10 pllCtrlSpiBusy R W I=i_pllCtrlSpiBusy_p
--   11:11 refDacSpiStart R W O=o_refDacSpiStart_p
--   12:12 refDacSpiBusy R W I=i_refDacSpiBusy_p
--   2:2 txGainSpiStart R W O=o_txGainSpiStart_p
--   3:3 txGainSpiBusy R I=i_txGainSpiBusy_p
--   31:13 rsvd2 R
--   6:4 RxGainSpiStart R W O=ov3_RxGainSpiStart_p
--   7:7 rxGainSpiBusy R W I=i_rxGainSpiBusy_p
--   9:8 pllCtrlSpiStart R W O=ov2_pllCtrlSpiStart_p

-- BASEADDR + 0x24   TXIQGAINIMBALANCE    Gain correction on I to fix IQ gain imbalance
--   12:0 IQGainImb R W O=ov13_IQGainImb_p
--   31:13 rsvd R

-- BASEADDR + 0x28   TXIQPHASEIMBALANCE    IQ phase constants to apply
--   12:0 IQPhaseImbCos R W O=ov13_IQPhaseImbCos_p
--   15:13 rsvd0 R
--   28:16 IQPhaseImbSin R W O=ov13_IQPhaseImbSin_p
--   31:29 rsvd1 R

-- BASEADDR + 0x2c   TXIQIMBALANCEBACKOFF    Backoff correction to not saturate value
--   12:0 IQImbBackOff R W O=ov13_IQImbBackOff_p
--   31:13 rsvd R

-- BASEADDR + 0x30   RSVD0    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x34   RSVD1    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x38   RXDCLEVEL    Give the RXI and RXQ DC level
--   11:0 RxIDcVal R I=iv12_RxIDcVal_p
--   15:12 rsvd0 R
--   27:16 RxQDcVal R I=iv12_RxQDcVal_p
--   31:28 rsvd1 R

-- BASEADDR + 0x3c   RXERF    Give the ERF as specified in the calibration guide of the LMS6002D
--   22:0 ERF R I=iv23_ERF_p
--   31:23 rsvd R

-- BASEADDR + 0x40   RSVD2    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x44   RSVD3    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x48   RSVD4    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x4c   RSVD5    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x50   RSVD6    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x54   RSVD7    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x58   RSVD8    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x5c   RSVD9    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x60   RSVD10    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x64   ERR_FCT_REG0    Error Function control
--   0:0 RXERRFCT_START R W O=o_RXERRFCT_START_p
--   1:1 RXERRFCT_DONE R I=i_RXERRFCT_DONE_p
--   15:3 rsvd R
--   2:2 RXERRFCT_FREQ_WEN R W O=o_RXERRFCT_FREQ_WEN_p
--   29:16 RXERRFCT_NB_POINT R W O=ov14_RXERRFCT_NB_POINT_p
--   31:30 rsvd R

-- BASEADDR + 0x68   ERR_FCT_REG1    DDS Frequency
--   23:0 RXERRFCT_FREQ R W O=ov24_RXERRFCT_FREQ_p
--   31:24 rsvd R

-- BASEADDR + 0x6c   ERR_FCT_REG2    Err_I
--   31:0 RXERRFCT_ERR_I R I=iv32_RXERRFCT_ERR_I_p

-- BASEADDR + 0x70   ERR_FCT_REG3    Err_Q
--   31:0 RXERRFCT_ERR_Q R I=iv32_RXERRFCT_ERR_Q_p

-- BASEADDR + 0x74   ADC_IDELAY_CTRL    Control ADC IDELAY values
--   31:10 rsvd0 R
--   4:0 AdcIdelayValue R W O=ov5_AdcIdelayValue_p
--   9:5 AdcClkIdelayValue R W O=ov5_AdcClkIdelayValue_p

-- BASEADDR + 0x78   RSVD12    Reserved
--   31:0 rsvd0 R

-- BASEADDR + 0x7c   RSVD13    Reserved
--   31:0 rsvd0 R

--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library proc_common_v3_00_a;
use proc_common_v3_00_a.proc_common_pkg.all;

-- DO NOT EDIT ABOVE THIS LINE --------------------

--USER libraries added here

------------------------------------------------------------------------------
-- Entity section
------------------------------------------------------------------------------
-- Definition of Generics:
--   C_NUM_REG                    -- Number of software accessible registers
--   C_SLV_DWIDTH                 -- Slave interface data bus width
--
-- Definition of Ports:
--   Bus2IP_Clk                   -- Bus to IP clock
--   Bus2IP_Resetn                -- Bus to IP reset
--   Bus2IP_Data                  -- Bus to IP data bus
--   Bus2IP_BE                    -- Bus to IP byte enables
--   Bus2IP_RdCE                  -- Bus to IP read chip enable
--   Bus2IP_WrCE                  -- Bus to IP write chip enable
--   IP2Bus_Data                  -- IP to Bus data bus
--   IP2Bus_RdAck                 -- IP to Bus read transfer acknowledgement
--   IP2Bus_WrAck                 -- IP to Bus write transfer acknowledgement
--   IP2Bus_Error                 -- IP to Bus error response
------------------------------------------------------------------------------

entity user_logic is
  generic
  (
    -- ADD USER GENERICS BELOW THIS LINE ---------------
    --USER generics added here
    -- ADD USER GENERICS ABOVE THIS LINE ---------------

    -- DO NOT EDIT BELOW THIS LINE ---------------------
    -- Bus protocol parameters, do not add to or delete
    C_NUM_REG                      : integer              := 32;
    C_SLV_DWIDTH                   : integer              := 32
    -- DO NOT EDIT ABOVE THIS LINE ---------------------
  );
  port
  (
    -- ADD USER PORTS BELOW THIS LINE ------------------
    --USER ports added here
    -- ADD USER PORTS ABOVE THIS LINE ------------------
    -- User ports
  i_CoreReset_p : in std_logic;

    o_TxEnable_p : out std_logic;
    o_RxEnable_p : out std_logic;
    ov2_ClkMuxSout_p : out std_logic_vector(1 downto 0);
    o_ClkMuxLoad_p : out std_logic;
    o_ClkMuxConfig_p : out std_logic;
    i_PLLLock_p : in std_logic;
    i_ovrAdcI_p : in std_logic;
    i_ovrAdcQ_p : in std_logic;
    i_ovrDacI_p : in std_logic;
    i_ovrDacQ_p : in std_logic;
    i_fmcPps_p : in std_logic;
    o_LimeReset_p : out std_logic;
    o_ResetOvr_p : out std_logic;
    o_DesignClkEn_p : out std_logic;
    o_CoreResetPulse_p : out std_logic;
    o_RstFifo_p : out std_logic;
    ov5_FpgaControl_p : out std_logic_vector(4 downto 0);
    ov2_ClkMuxSin_p : out std_logic_vector(1 downto 0);
    ov24_ddsfreq_p : out std_logic_vector(23 downto 0);
    ov3_dacOutSel_p : out std_logic_vector(2 downto 0);
    ov16_limeSpiDataIn_p : out std_logic_vector(15 downto 0);
    iv16_limeSpiDataOut_p : in std_logic_vector(15 downto 0);
    ov6_txGainSpiData_p : out std_logic_vector(5 downto 0);
    ov6_rxGainSpiData_p : out std_logic_vector(5 downto 0);
    ov32_pllCtrlSpiDataIn_p : out std_logic_vector(31 downto 0);
    iv32_pllCtrlSpiDataOut_p : in std_logic_vector(31 downto 0);
    ov16_refDacSpiData_p : out std_logic_vector(15 downto 0);
    iv16_refDacSpiData_p : in std_logic_vector(15 downto 0);
    o_limeSpiStart_p : out std_logic;
    i_limeSpiBusy_p : in std_logic;
    i_pllCtrlSpiBusy_p : in std_logic;
    o_refDacSpiStart_p : out std_logic;
    i_refDacSpiBusy_p : in std_logic;
    o_txGainSpiStart_p : out std_logic;
    i_txGainSpiBusy_p : in std_logic;
    ov3_RxGainSpiStart_p : out std_logic_vector(2 downto 0);
    i_rxGainSpiBusy_p : in std_logic;
    ov2_pllCtrlSpiStart_p : out std_logic_vector(1 downto 0);
    ov13_IQGainImb_p : out std_logic_vector(12 downto 0);
    ov13_IQPhaseImbCos_p : out std_logic_vector(12 downto 0);
    ov13_IQPhaseImbSin_p : out std_logic_vector(12 downto 0);
    ov13_IQImbBackOff_p : out std_logic_vector(12 downto 0);
    iv12_RxIDcVal_p : in std_logic_vector(11 downto 0);
    iv12_RxQDcVal_p : in std_logic_vector(11 downto 0);
    iv23_ERF_p : in std_logic_vector(22 downto 0);
    o_RXERRFCT_START_p : out std_logic;
    i_RXERRFCT_DONE_p : in std_logic;
    o_RXERRFCT_FREQ_WEN_p : out std_logic;
    ov14_RXERRFCT_NB_POINT_p : out std_logic_vector(13 downto 0);
    ov24_RXERRFCT_FREQ_p : out std_logic_vector(23 downto 0);
    iv32_RXERRFCT_ERR_I_p : in std_logic_vector(31 downto 0);
    iv32_RXERRFCT_ERR_Q_p : in std_logic_vector(31 downto 0);
    ov5_AdcIdelayValue_p : out std_logic_vector(4 downto 0);
    ov5_AdcClkIdelayValue_p : out std_logic_vector(4 downto 0);
    -- Bus protocol ports, do not add to or delete
    Bus2IP_Clk                     : in  std_logic;
    Bus2IP_Resetn                  : in  std_logic;
    Bus2IP_Data                    : in  std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    Bus2IP_BE                      : in  std_logic_vector(C_SLV_DWIDTH/8-1 downto 0);
    Bus2IP_RdCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    Bus2IP_WrCE                    : in  std_logic_vector(C_NUM_REG-1 downto 0);
    IP2Bus_Data                    : out std_logic_vector(C_SLV_DWIDTH-1 downto 0);
    IP2Bus_RdAck                   : out std_logic;
    IP2Bus_WrAck                   : out std_logic;
    IP2Bus_Error                   : out std_logic
  );

 attribute MAX_FANOUT : string;
 attribute SIGIS : string;
 attribute SIGIS of Bus2IP_Clk    : signal is "CLK";
 attribute SIGIS of Bus2IP_Resetn : signal is "RST";

end entity user_logic;

------------------------------------------------------------------------------
-- Architecture section
------------------------------------------------------------------------------

architecture IMP of user_logic is

-------------------------------------------------------------------------------
-- Constant declarations
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
--     ************** Function declaratin *******************                   
-- Return a std_logic_vector with only one bit set to one.
-- The argument BitPosition represent the bit position to set to one, starting with 0.
-- The argument Width represent the width of the returned std_logic_vector.
-------------------------------------------------------------------------------
  function OneHotVector( BitPosition : integer;                              
                Width : integer)                                             
                return std_logic_vector                                      
  is                                                                         
    variable Result                   : std_logic_vector(Width - 1 downto 0);

  begin                        
    Result := (others => '0'); 
    Result(BitPosition) := '1';
    return Result;             
  end OneHotVector;            
-------------------------------------------------------------------------------
-- Signal and Type Declarations
-------------------------------------------------------------------------------

  signal TxEnable_s                     : std_logic;
  signal RxEnable_s                     : std_logic;
  signal v2_ClkMuxSout_s                     : std_logic_vector(1 downto 0);
  signal ClkMuxLoad_s                     : std_logic;
  signal ClkMuxConfig_s                     : std_logic;
  signal LimeReset_s                     : std_logic;
  signal ResetOvr_s                     : std_logic;
  signal DesignClkEn_s                     : std_logic;
  signal CoreResetPulse_s                     : std_logic;
  signal RstFifo_s                     : std_logic;
  signal v5_FpgaControl_s                     : std_logic_vector(4 downto 0);
  signal v2_ClkMuxSin_s                     : std_logic_vector(1 downto 0);
  signal v24_ddsfreq_s                     : std_logic_vector(23 downto 0);
  signal v3_dacOutSel_s                     : std_logic_vector(2 downto 0);
  signal v16_limeSpiDataIn_s                     : std_logic_vector(15 downto 0);
  signal v6_txGainSpiData_s                     : std_logic_vector(5 downto 0);
  signal v6_rxGainSpiData_s                     : std_logic_vector(5 downto 0);
  signal v32_pllCtrlSpiDataIn_s                     : std_logic_vector(31 downto 0);
  signal v16_refDacSpiData_s                     : std_logic_vector(15 downto 0);
  signal limeSpiStart_s                     : std_logic;
  signal pllCtrlSpiBusy_s                     : std_logic;
  signal refDacSpiStart_s                     : std_logic;
  signal refDacSpiBusy_s                     : std_logic;
  signal txGainSpiStart_s                     : std_logic;
  signal v3_RxGainSpiStart_s                     : std_logic_vector(2 downto 0);
  signal rxGainSpiBusy_s                     : std_logic;
  signal v2_pllCtrlSpiStart_s                     : std_logic_vector(1 downto 0);
  signal v13_IQGainImb_s                     : std_logic_vector(12 downto 0);
  signal v13_IQPhaseImbCos_s                     : std_logic_vector(12 downto 0);
  signal v13_IQPhaseImbSin_s                     : std_logic_vector(12 downto 0);
  signal v13_IQImbBackOff_s                     : std_logic_vector(12 downto 0);
  signal RXERRFCT_START_s                     : std_logic;
  signal RXERRFCT_FREQ_WEN_s                     : std_logic;
  signal v14_RXERRFCT_NB_POINT_s                     : std_logic_vector(13 downto 0);
  signal v24_RXERRFCT_FREQ_s                     : std_logic_vector(23 downto 0);
  signal v5_AdcIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal v5_AdcClkIdelayValue_s                     : std_logic_vector(4 downto 0);
  signal slv_reg_write_sel              : std_logic_vector(31 downto 0);
  signal slv_reg_read_sel               : std_logic_vector(31 downto 0);
  signal slv_ip2bus_data                : std_logic_vector(C_SLV_DWIDTH-1 downto 0);
  signal slv_read_ack                   : std_logic;
  signal slv_write_ack                  : std_logic;

------------------------------------------------------------------------------
begin
------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Begin architecture
-------------------------------------------------------------------------------

-- swap bits
WrCeBitSwap: for i in 0 to slv_reg_write_sel'high generate
  slv_reg_write_sel(i) <= Bus2IP_WrCE(slv_reg_write_sel'high - i);
end generate WrCeBitSwap;

RdCeBitSwap: for i in 0 to slv_reg_read_sel'high generate
  slv_reg_read_sel(i)  <= Bus2IP_RdCE(slv_reg_read_sel'high - i);
end generate RdCeBitSwap;

-- generate write/read ack
  slv_write_ack <=   Bus2IP_WrCE(0) or   Bus2IP_WrCE(1) or   Bus2IP_WrCE(2) or   Bus2IP_WrCE(3) or   Bus2IP_WrCE(4) or   Bus2IP_WrCE(5) or   Bus2IP_WrCE(6) or   Bus2IP_WrCE(7) or   Bus2IP_WrCE(8) or   Bus2IP_WrCE(9) or   Bus2IP_WrCE(10) or   Bus2IP_WrCE(11) or   Bus2IP_WrCE(12) or   Bus2IP_WrCE(13) or   Bus2IP_WrCE(14) or   Bus2IP_WrCE(15) or   Bus2IP_WrCE(16) or   Bus2IP_WrCE(17) or   Bus2IP_WrCE(18) or   Bus2IP_WrCE(19) or   Bus2IP_WrCE(20) or   Bus2IP_WrCE(21) or   Bus2IP_WrCE(22) or   Bus2IP_WrCE(23) or   Bus2IP_WrCE(24) or   Bus2IP_WrCE(25) or   Bus2IP_WrCE(26) or   Bus2IP_WrCE(27) or   Bus2IP_WrCE(28) or   Bus2IP_WrCE(29) or   Bus2IP_WrCE(30) or   Bus2IP_WrCE(31);
  slv_read_ack  <=   Bus2IP_RdCE(0) or   Bus2IP_RdCE(1) or   Bus2IP_RdCE(2) or   Bus2IP_RdCE(3) or   Bus2IP_RdCE(4) or   Bus2IP_RdCE(5) or   Bus2IP_RdCE(6) or   Bus2IP_RdCE(7) or   Bus2IP_RdCE(8) or   Bus2IP_RdCE(9) or   Bus2IP_RdCE(10) or   Bus2IP_RdCE(11) or   Bus2IP_RdCE(12) or   Bus2IP_RdCE(13) or   Bus2IP_RdCE(14) or   Bus2IP_RdCE(15) or   Bus2IP_RdCE(16) or   Bus2IP_RdCE(17) or   Bus2IP_RdCE(18) or   Bus2IP_RdCE(19) or   Bus2IP_RdCE(20) or   Bus2IP_RdCE(21) or   Bus2IP_RdCE(22) or   Bus2IP_RdCE(23) or   Bus2IP_RdCE(24) or   Bus2IP_RdCE(25) or   Bus2IP_RdCE(26) or   Bus2IP_RdCE(27) or   Bus2IP_RdCE(28) or   Bus2IP_RdCE(29) or   Bus2IP_RdCE(30) or   Bus2IP_RdCE(31);

 -- implement slave model software accessible register(s)
 SLAVE_REG_WRITE_PROC : process( Bus2IP_Clk ) is
 begin

  if Bus2IP_Clk'event and Bus2IP_Clk = '1' then
    if Bus2IP_Resetn = '0' then
      TxEnable_s <= '0';
      RxEnable_s <= '0';
      v2_ClkMuxSout_s <=  "00";
      ClkMuxLoad_s <=  '0';
      ClkMuxConfig_s <=  '0';
      LimeReset_s <= '0';
      ResetOvr_s <=  '0';
      DesignClkEn_s <=  '0';
      CoreResetPulse_s <= '0';
      RstFifo_s <=  '1';
      v5_FpgaControl_s <= "00000";
      v2_ClkMuxSin_s <= "00";
      v24_ddsfreq_s <= X"000000";
      v3_dacOutSel_s <= "000";
      v16_limeSpiDataIn_s <= X"0000";
      v6_txGainSpiData_s <= "000000";
      v6_rxGainSpiData_s <= "000000";
      v32_pllCtrlSpiDataIn_s <= X"00000000";
      v16_refDacSpiData_s <= X"0000";
      limeSpiStart_s <= '0';
--      pllCtrlSpiBusy_s <= '0';
      refDacSpiStart_s <= '0';
--      refDacSpiBusy_s <= '0';
      txGainSpiStart_s <= '0';
      v3_RxGainSpiStart_s <= "000";
--      rxGainSpiBusy_s <= '0';
      v2_pllCtrlSpiStart_s <= "00";
      v13_IQGainImb_s <= '0'& X"800";
      v13_IQPhaseImbCos_s <= '0'& X"800";
      v13_IQPhaseImbSin_s <= '0' & X"000";
      v13_IQImbBackOff_s <= '0' & X"800";
      RXERRFCT_START_s <= '0';
      RXERRFCT_FREQ_WEN_s <= '0';
      v14_RXERRFCT_NB_POINT_s <=  "00000000000000";
      v24_RXERRFCT_FREQ_s <= x"000000";
      v5_AdcIdelayValue_s <=  "00000";
      v5_AdcClkIdelayValue_s <=  "00000";

    else

  -- Synchronous reset
  if ( i_CoreReset_p = '1' ) then
    TxEnable_s <= '0';
    RxEnable_s <= '0';
    v2_ClkMuxSout_s <=  "00";
    ClkMuxLoad_s <=  '0';
    ClkMuxConfig_s <=  '0';
    LimeReset_s <= '0';
    ResetOvr_s <=  '0';
    DesignClkEn_s <=  '0';
    CoreResetPulse_s <= '0';
    RstFifo_s <=  '1';
    v5_FpgaControl_s <= "00000";
    v2_ClkMuxSin_s <= "00";
    v24_ddsfreq_s <= X"000000";
    v3_dacOutSel_s <= "000";
    v16_limeSpiDataIn_s <= X"0000";
    v6_txGainSpiData_s <= "000000";
    v6_rxGainSpiData_s <= "000000";
    v32_pllCtrlSpiDataIn_s <= X"00000000";
    v16_refDacSpiData_s <= X"0000";
    limeSpiStart_s <= '0';
--    pllCtrlSpiBusy_s <= '0';
    refDacSpiStart_s <= '0';
--    refDacSpiBusy_s <= '0';
    txGainSpiStart_s <= '0';
    v3_RxGainSpiStart_s <= "000";
--    rxGainSpiBusy_s <= '0';
    v2_pllCtrlSpiStart_s <= "00";
    v13_IQGainImb_s <= '0'& X"800";
    v13_IQPhaseImbCos_s <= '0'& X"800";
    v13_IQPhaseImbSin_s <= '0' & X"000";
    v13_IQImbBackOff_s <= '0' & X"800";
    RXERRFCT_START_s <= '0';
    RXERRFCT_FREQ_WEN_s <= '0';
    v14_RXERRFCT_NB_POINT_s <=  "00000000000000";
    v24_RXERRFCT_FREQ_s <= x"000000";
    v5_AdcIdelayValue_s <=  "00000";
    v5_AdcClkIdelayValue_s <=  "00000";
  end if;

  CoreResetPulse_s <= '0';
      case slv_reg_write_sel is

        when OneHotVector(1,32) =>
          if (Bus2IP_BE(0) = '1') then
            TxEnable_s <= Bus2IP_Data(0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            RxEnable_s <= Bus2IP_Data(1);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v2_ClkMuxSout_s <= Bus2IP_Data(11 downto 10);
          end if;
          if (Bus2IP_BE(1) = '1') then
            ClkMuxLoad_s <= Bus2IP_Data(12);
          end if;
          if (Bus2IP_BE(1) = '1') then
            ClkMuxConfig_s <= Bus2IP_Data(13);
          end if;
          if (Bus2IP_BE(0) = '1') then
            LimeReset_s <= Bus2IP_Data(2);
          end if;
          if (Bus2IP_BE(2) = '1') then
            ResetOvr_s <= Bus2IP_Data(20);
          end if;
          if (Bus2IP_BE(3) = '1') then
            DesignClkEn_s <= Bus2IP_Data(25);
          end if;
          if (Bus2IP_BE(3) = '1') then
            CoreResetPulse_s <= Bus2IP_Data(26);
          end if;
          if (Bus2IP_BE(3) = '1') then
            RstFifo_s <= Bus2IP_Data(27);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v5_FpgaControl_s <= Bus2IP_Data(7 downto 3);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v2_ClkMuxSin_s <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(2,32) =>
          if (Bus2IP_BE(0) = '1') then
            v24_ddsfreq_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v24_ddsfreq_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v24_ddsfreq_s(23 downto 16) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v3_dacOutSel_s <= Bus2IP_Data(26 downto 24);
          end if;

        when OneHotVector(3,32) =>
          if (Bus2IP_BE(0) = '1') then
            v16_limeSpiDataIn_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v16_limeSpiDataIn_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;

        when OneHotVector(4,32) =>
          if (Bus2IP_BE(0) = '1') then
            v6_txGainSpiData_s <= Bus2IP_Data(5 downto 0);
          end if;

        when OneHotVector(5,32) =>
          if (Bus2IP_BE(0) = '1') then
            v6_rxGainSpiData_s <= Bus2IP_Data(5 downto 0);
          end if;

        when OneHotVector(6,32) =>
          if (Bus2IP_BE(0) = '1') then
            v32_pllCtrlSpiDataIn_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v32_pllCtrlSpiDataIn_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v32_pllCtrlSpiDataIn_s(23 downto 16) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v32_pllCtrlSpiDataIn_s(31 downto 24) <= Bus2IP_Data(31 downto 24);
          end if;

        when OneHotVector(7,32) =>
          if (Bus2IP_BE(0) = '1') then
            v16_refDacSpiData_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v16_refDacSpiData_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;

        when OneHotVector(8,32) =>
          if (Bus2IP_BE(0) = '1') then
            limeSpiStart_s <= Bus2IP_Data(0);
          end if;
          if (Bus2IP_BE(1) = '1') then
--            pllCtrlSpiBusy_s <= Bus2IP_Data(10);
          end if;
          if (Bus2IP_BE(1) = '1') then
            refDacSpiStart_s <= Bus2IP_Data(11);
          end if;
          if (Bus2IP_BE(1) = '1') then
--            refDacSpiBusy_s <= Bus2IP_Data(12);
          end if;
          if (Bus2IP_BE(0) = '1') then
            txGainSpiStart_s <= Bus2IP_Data(2);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v3_RxGainSpiStart_s <= Bus2IP_Data(6 downto 4);
          end if;
          if (Bus2IP_BE(0) = '1') then
--            rxGainSpiBusy_s <= Bus2IP_Data(7);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v2_pllCtrlSpiStart_s <= Bus2IP_Data(9 downto 8);
          end if;

        when OneHotVector(9,32) =>
          if (Bus2IP_BE(0) = '1') then
            v13_IQGainImb_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v13_IQGainImb_s(12 downto 8) <= Bus2IP_Data(12 downto 8);
          end if;

        when OneHotVector(10,32) =>
          if (Bus2IP_BE(0) = '1') then
            v13_IQPhaseImbCos_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v13_IQPhaseImbCos_s(12 downto 8) <= Bus2IP_Data(12 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v13_IQPhaseImbSin_s(7 downto 0) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v13_IQPhaseImbSin_s(12 downto 8) <= Bus2IP_Data(28 downto 24);
          end if;

        when OneHotVector(11,32) =>
          if (Bus2IP_BE(0) = '1') then
            v13_IQImbBackOff_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v13_IQImbBackOff_s(12 downto 8) <= Bus2IP_Data(12 downto 8);
          end if;

        when OneHotVector(25,32) =>
          if (Bus2IP_BE(0) = '1') then
            RXERRFCT_START_s <= Bus2IP_Data(0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            RXERRFCT_FREQ_WEN_s <= Bus2IP_Data(2);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v14_RXERRFCT_NB_POINT_s(7 downto 0) <= Bus2IP_Data(23 downto 16);
          end if;
          if (Bus2IP_BE(3) = '1') then
            v14_RXERRFCT_NB_POINT_s(13 downto 8) <= Bus2IP_Data(29 downto 24);
          end if;

        when OneHotVector(26,32) =>
          if (Bus2IP_BE(0) = '1') then
            v24_RXERRFCT_FREQ_s(7 downto 0) <= Bus2IP_Data(7 downto 0);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v24_RXERRFCT_FREQ_s(15 downto 8) <= Bus2IP_Data(15 downto 8);
          end if;
          if (Bus2IP_BE(2) = '1') then
            v24_RXERRFCT_FREQ_s(23 downto 16) <= Bus2IP_Data(23 downto 16);
          end if;

        when OneHotVector(29,32) =>
          if (Bus2IP_BE(0) = '1') then
            v5_AdcIdelayValue_s <= Bus2IP_Data(4 downto 0);
          end if;
          if (Bus2IP_BE(0) = '1') then
            v5_AdcClkIdelayValue_s(2 downto 0) <= Bus2IP_Data(7 downto 5);
          end if;
          if (Bus2IP_BE(1) = '1') then
            v5_AdcClkIdelayValue_s(4 downto 3) <= Bus2IP_Data(9 downto 8);
          end if;
        when others =>
          null;
      end case;
    end if;
  end if;

 end process SLAVE_REG_WRITE_PROC;

 -- implement slave model software accessible register(s) read mux
SLAVE_REG_READ_PROC : process( slv_reg_read_sel, TxEnable_s, RxEnable_s, v2_ClkMuxSout_s, ClkMuxLoad_s, ClkMuxConfig_s, i_PLLLock_p, i_ovrAdcI_p, i_ovrAdcQ_p, i_ovrDacI_p, i_ovrDacQ_p, i_fmcPps_p, LimeReset_s, ResetOvr_s, DesignClkEn_s, RstFifo_s, v5_FpgaControl_s, v2_ClkMuxSin_s, v24_ddsfreq_s, v3_dacOutSel_s, iv16_limeSpiDataOut_p, v6_txGainSpiData_s, v6_rxGainSpiData_s, iv32_pllCtrlSpiDataOut_p, limeSpiStart_s, i_limeSpiBusy_p, i_pllCtrlSpiBusy_p, refDacSpiStart_s, i_refDacSpiBusy_p, txGainSpiStart_s, i_txGainSpiBusy_p, v3_RxGainSpiStart_s, i_rxGainSpiBusy_p, v2_pllCtrlSpiStart_s, v13_IQGainImb_s, v13_IQPhaseImbCos_s, v13_IQPhaseImbSin_s, v13_IQImbBackOff_s, iv12_RxIDcVal_p, RXERRFCT_START_s, i_RXERRFCT_DONE_p, RXERRFCT_FREQ_WEN_s, v14_RXERRFCT_NB_POINT_s, v24_RXERRFCT_FREQ_s, iv32_RXERRFCT_ERR_I_p, iv32_RXERRFCT_ERR_Q_p, iv16_refDacSpiData_p, v5_AdcIdelayValue_s, v5_AdcClkIdelayValue_s) is
 begin
   case slv_reg_read_sel is

        when OneHotVector(0,32) =>
          slv_ip2bus_data(31 downto 0) <= X"FCC10200";

        when OneHotVector(1,32) =>
          slv_ip2bus_data(0) <= TxEnable_s;
          slv_ip2bus_data(1) <= RxEnable_s;
          slv_ip2bus_data(11 downto 10) <= v2_ClkMuxSout_s;
          slv_ip2bus_data(12) <= ClkMuxLoad_s;
          slv_ip2bus_data(13) <= ClkMuxConfig_s;
          slv_ip2bus_data(14) <= i_PLLLock_p;
          slv_ip2bus_data(15) <= i_ovrAdcI_p;
          slv_ip2bus_data(16) <= i_ovrAdcQ_p;
          slv_ip2bus_data(17) <= i_ovrDacI_p;
          slv_ip2bus_data(18) <= i_ovrDacQ_p;
          slv_ip2bus_data(19) <= i_fmcPps_p;
          slv_ip2bus_data(2) <= LimeReset_s;
          slv_ip2bus_data(20) <= ResetOvr_s;
          slv_ip2bus_data(24 downto 21) <= "0000";
          slv_ip2bus_data(25) <= DesignClkEn_s;
          slv_ip2bus_data(27) <= RstFifo_s;
          slv_ip2bus_data(31 downto 28) <= "0000";
          slv_ip2bus_data(7 downto 3) <= v5_FpgaControl_s;
          slv_ip2bus_data(9 downto 8) <= v2_ClkMuxSin_s;

        when OneHotVector(2,32) =>
          slv_ip2bus_data(23 downto 0) <= v24_ddsfreq_s;
          slv_ip2bus_data(26 downto 24) <= v3_dacOutSel_s;
          slv_ip2bus_data(31 downto 27) <= "00000";

        when OneHotVector(3,32) =>
          slv_ip2bus_data(15 downto 0) <= iv16_limeSpiDataOut_p;
          slv_ip2bus_data(31 downto 16) <= X"0000";

        when OneHotVector(4,32) =>
          slv_ip2bus_data(31 downto 6) <= X"0000" & "0000000000";
          slv_ip2bus_data(5 downto 0) <= v6_txGainSpiData_s;

        when OneHotVector(5,32) =>
          slv_ip2bus_data(31 downto 6) <= X"0000" & "0000000000";
          slv_ip2bus_data(5 downto 0) <= v6_rxGainSpiData_s;

        when OneHotVector(6,32) =>
          slv_ip2bus_data(31 downto 0) <= iv32_pllCtrlSpiDataOut_p;

        when OneHotVector(7,32) =>
          slv_ip2bus_data(15 downto 0) <= iv16_refDacSpiData_p;
          slv_ip2bus_data(31 downto 16) <= X"0000";

        when OneHotVector(8,32) =>
          slv_ip2bus_data(0) <= limeSpiStart_s;
          slv_ip2bus_data(1) <= i_limeSpiBusy_p;
          slv_ip2bus_data(10) <= i_pllCtrlSpiBusy_p;
          slv_ip2bus_data(11) <= refDacSpiStart_s;
          slv_ip2bus_data(12) <= i_refDacSpiBusy_p;
          slv_ip2bus_data(2) <= txGainSpiStart_s;
          slv_ip2bus_data(3) <= i_txGainSpiBusy_p;
          slv_ip2bus_data(31 downto 13) <= "0000000000000000000";
          slv_ip2bus_data(6 downto 4) <= v3_RxGainSpiStart_s;
          slv_ip2bus_data(7) <= i_rxGainSpiBusy_p;
          slv_ip2bus_data(9 downto 8) <= v2_pllCtrlSpiStart_s;

        when OneHotVector(9,32) =>
          slv_ip2bus_data(12 downto 0) <= v13_IQGainImb_s;
          slv_ip2bus_data(31 downto 13) <= X"0000" & "000";

        when OneHotVector(10,32) =>
          slv_ip2bus_data(12 downto 0) <= v13_IQPhaseImbCos_s;
          slv_ip2bus_data(15 downto 13) <= "000";
          slv_ip2bus_data(28 downto 16) <= v13_IQPhaseImbSin_s;
          slv_ip2bus_data(31 downto 29) <= "000";

        when OneHotVector(11,32) =>
          slv_ip2bus_data(12 downto 0) <= v13_IQImbBackOff_s;
          slv_ip2bus_data(31 downto 13) <= X"0000" & "000";

        when OneHotVector(12,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(13,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(14,32) =>
          slv_ip2bus_data(11 downto 0) <= iv12_RxIDcVal_p;
          slv_ip2bus_data(15 downto 12) <=  X"0";
          slv_ip2bus_data(27 downto 16) <= iv12_RxQDcVal_p;
          slv_ip2bus_data(31 downto 28) <= X"0";

        when OneHotVector(15,32) =>
          slv_ip2bus_data(22 downto 0) <= iv23_ERF_p;
          slv_ip2bus_data(31 downto 23) <= "000000000";

        when OneHotVector(16,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(17,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(18,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(19,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(20,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(21,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(22,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(23,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(24,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(25,32) =>
          slv_ip2bus_data(0) <= RXERRFCT_START_s;
          slv_ip2bus_data(1) <= i_RXERRFCT_DONE_p;
          slv_ip2bus_data(15 downto 3) <=  "0000000000000";
          slv_ip2bus_data(2) <= RXERRFCT_FREQ_WEN_s;
          slv_ip2bus_data(29 downto 16) <= v14_RXERRFCT_NB_POINT_s;
          slv_ip2bus_data(31 downto 30) <=  "00";

        when OneHotVector(26,32) =>
          slv_ip2bus_data(23 downto 0) <= v24_RXERRFCT_FREQ_s;
          slv_ip2bus_data(31 downto 24) <=  X"00";

        when OneHotVector(27,32) =>
          slv_ip2bus_data(31 downto 0) <= iv32_RXERRFCT_ERR_I_p;

        when OneHotVector(28,32) =>
          slv_ip2bus_data(31 downto 0) <= iv32_RXERRFCT_ERR_Q_p;

        when OneHotVector(29,32) =>
          slv_ip2bus_data(31 downto 10) <=  "0000000000000000000000";
          slv_ip2bus_data(4 downto 0) <= v5_AdcIdelayValue_s;
          slv_ip2bus_data(9 downto 5) <= v5_AdcClkIdelayValue_s;

        when OneHotVector(30,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";

        when OneHotVector(31,32) =>
          slv_ip2bus_data(31 downto 0) <=  X"00000000";
        when others =>
          slv_ip2bus_data <= (others => '0');
      end case;

 end process SLAVE_REG_READ_PROC;

------------------------------------------
-- drive IP to Bus signals
------------------------------------------
IP2Bus_Data  <= slv_ip2bus_data when slv_read_ack = '1' else (others => '0');
IP2Bus_WrAck <= slv_write_ack;
IP2Bus_RdAck <= slv_read_ack;
IP2Bus_Error <= '0';

------------------------------------------
-- Output assignments
------------------------------------------
o_TxEnable_p <= TxEnable_s;
o_RxEnable_p <= RxEnable_s;
ov2_ClkMuxSout_p <= v2_ClkMuxSout_s;
o_ClkMuxLoad_p <= ClkMuxLoad_s;
o_ClkMuxConfig_p <= ClkMuxConfig_s;
o_LimeReset_p <= LimeReset_s;
o_ResetOvr_p <= ResetOvr_s;
o_DesignClkEn_p <= DesignClkEn_s;
o_CoreResetPulse_p <= CoreResetPulse_s;
o_RstFifo_p <= RstFifo_s;
ov5_FpgaControl_p <= v5_FpgaControl_s;
ov2_ClkMuxSin_p <= v2_ClkMuxSin_s;
ov24_ddsfreq_p <= v24_ddsfreq_s;
ov3_dacOutSel_p <= v3_dacOutSel_s;
ov16_limeSpiDataIn_p <= v16_limeSpiDataIn_s;
ov6_txGainSpiData_p <= v6_txGainSpiData_s;
ov6_rxGainSpiData_p <= v6_rxGainSpiData_s;
ov32_pllCtrlSpiDataIn_p <= v32_pllCtrlSpiDataIn_s;
ov16_refDacSpiData_p <= v16_refDacSpiData_s;
o_limeSpiStart_p <= limeSpiStart_s;
o_refDacSpiStart_p <= refDacSpiStart_s;
o_txGainSpiStart_p <= txGainSpiStart_s;
ov3_RxGainSpiStart_p <= v3_RxGainSpiStart_s;
ov2_pllCtrlSpiStart_p <= v2_pllCtrlSpiStart_s;
ov13_IQGainImb_p <= v13_IQGainImb_s;
ov13_IQPhaseImbCos_p <= v13_IQPhaseImbCos_s;
ov13_IQPhaseImbSin_p <= v13_IQPhaseImbSin_s;
ov13_IQImbBackOff_p <= v13_IQImbBackOff_s;
o_RXERRFCT_START_p <= RXERRFCT_START_s;
o_RXERRFCT_FREQ_WEN_p <= RXERRFCT_FREQ_WEN_s;
ov14_RXERRFCT_NB_POINT_p <= v14_RXERRFCT_NB_POINT_s;
ov24_RXERRFCT_FREQ_p <= v24_RXERRFCT_FREQ_s;
ov5_AdcIdelayValue_p <= v5_AdcIdelayValue_s;
ov5_AdcClkIdelayValue_p <= v5_AdcClkIdelayValue_s;

end IMP;

