-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.5
--  \   \         Application :  Virtex-6 FPGA GTX Transceiver Wizard
--  /   /         Filename : gtx_wrapper.vhd
-- /___/   /\     Timestamp :
-- \   \  /  \
--  \___\/\___\
--
--
-- Module GTX_WRAPPER (a GTX Wrapper)
-- Generated by Xilinx Virtex-6 FPGA GTX Transceiver Wizard
-- 
-- 
-- (c) Copyright 2009 - 2010 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity GTX_WRAPPER is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0 -- Set to 1 to speed up sim reset
);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX0  (X0Y0)

    ------------------------ Loopback and Powerdown Ports ----------------------
    GTX0_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    GTX0_RXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    GTX0_TXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GTX0_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GTX0_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    GTX0_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GTX0_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GTX0_RXCHANBONDSEQ_OUT                  : out  std_logic;
    GTX0_RXCHBONDI_IN                       : in   std_logic_vector(3 downto 0);
    GTX0_RXCHBONDLEVEL_IN                   : in   std_logic_vector(2 downto 0);
    GTX0_RXCHBONDMASTER_IN                  : in   std_logic;
    GTX0_RXCHBONDO_OUT                      : out  std_logic_vector(3 downto 0);
    GTX0_RXCHBONDSLAVE_IN                   : in   std_logic;
    GTX0_RXENCHANSYNC_IN                    : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GTX0_RXCLKCORCNT_OUT                    : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------    
    GTX0_RXBYTEISALIGNED_OUT                : out  std_logic;
    GTX0_RXBYTEREALIGN_OUT                  : out  std_logic;
    GTX0_RXCOMMADET_OUT                     : out  std_logic;
    GTX0_RXENMCOMMAALIGN_IN                 : in   std_logic;
    GTX0_RXENPCOMMAALIGN_IN                 : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GTX0_PRBSCNTRESET_IN                    : in   std_logic;
    GTX0_RXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX0_RXPRBSERR_OUT                      : out  std_logic;    
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTX0_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    GTX0_RXRESET_IN                         : in   std_logic;
    GTX0_RXUSRCLK2_IN                       : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX0_RXCDRRESET_IN                      : in   std_logic;
    GTX0_RXELECIDLE_OUT                     : out  std_logic;
    GTX0_RXEQMIX_IN                         : in   std_logic_vector(2 downto 0);
    GTX0_RXN_IN                             : in   std_logic;
    GTX0_RXP_IN                             : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GTX0_RXBUFRESET_IN                      : in   std_logic;
    GTX0_RXBUFSTATUS_OUT                    : out  std_logic_vector(2 downto 0);
    GTX0_RXCHANISALIGNED_OUT                : out  std_logic;
    GTX0_RXCHANREALIGN_OUT                  : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    GTX0_RXLOSSOFSYNC_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTX0_GTXRXRESET_IN                      : in   std_logic;
    GTX0_MGTREFCLKRX_IN                     : in   std_logic;
    GTX0_PLLRXRESET_IN                      : in   std_logic;
    GTX0_RXPLLLKDET_OUT                     : out  std_logic;
    GTX0_RXRESETDONE_OUT                    : out  std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    GTX0_DADDR_IN                           : in   std_logic_vector(7 downto 0);
    GTX0_DCLK_IN                            : in   std_logic;
    GTX0_DEN_IN                             : in   std_logic;
    GTX0_DI_IN                              : in   std_logic_vector(15 downto 0);
    GTX0_DRDY_OUT                           : out  std_logic;
    GTX0_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GTX0_DWE_IN                             : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX0_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX0_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    GTX0_TXOUTCLK_OUT                       : out  std_logic;
    GTX0_TXRESET_IN                         : in   std_logic;
    GTX0_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX0_TXDIFFCTRL_IN                      : in   std_logic_vector(3 downto 0);
    GTX0_TXN_OUT                            : out  std_logic;
    GTX0_TXP_OUT                            : out  std_logic;
    GTX0_TXPOSTEMPHASIS_IN                  : in   std_logic_vector(4 downto 0);
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    GTX0_TXPREEMPHASIS_IN                   : in   std_logic_vector(3 downto 0);
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    GTX0_TXDLYALIGNDISABLE_IN               : in   std_logic;
    GTX0_TXDLYALIGNMONENB_IN                : in   std_logic;
    GTX0_TXDLYALIGNMONITOR_OUT              : out  std_logic_vector(7 downto 0);
    GTX0_TXDLYALIGNRESET_IN                 : in   std_logic;
    GTX0_TXENPMAPHASEALIGN_IN               : in   std_logic;
    GTX0_TXPMASETPHASE_IN                   : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX0_GTXTXRESET_IN                      : in   std_logic;
    GTX0_TXRESETDONE_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GTX0_TXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX0_TXPRBSFORCEERR_IN                  : in   std_logic;    
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GTX0_TXELECIDLE_IN                      : in   std_logic;



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX1  (X0Y1)

    ------------------------ Loopback and Powerdown Ports ----------------------
    GTX1_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    GTX1_RXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    GTX1_TXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GTX1_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GTX1_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    GTX1_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GTX1_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GTX1_RXCHANBONDSEQ_OUT                  : out  std_logic;
    GTX1_RXCHBONDI_IN                       : in   std_logic_vector(3 downto 0);
    GTX1_RXCHBONDLEVEL_IN                   : in   std_logic_vector(2 downto 0);
    GTX1_RXCHBONDMASTER_IN                  : in   std_logic;
    GTX1_RXCHBONDO_OUT                      : out  std_logic_vector(3 downto 0);
    GTX1_RXCHBONDSLAVE_IN                   : in   std_logic;
    GTX1_RXENCHANSYNC_IN                    : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GTX1_RXCLKCORCNT_OUT                    : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GTX1_RXBYTEISALIGNED_OUT                : out  std_logic;
    GTX1_RXBYTEREALIGN_OUT                  : out  std_logic;
    GTX1_RXCOMMADET_OUT                     : out  std_logic;
    GTX1_RXENMCOMMAALIGN_IN                 : in   std_logic;
    GTX1_RXENPCOMMAALIGN_IN                 : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GTX1_PRBSCNTRESET_IN                    : in   std_logic;
    GTX1_RXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX1_RXPRBSERR_OUT                      : out  std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTX1_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    GTX1_RXRESET_IN                         : in   std_logic;
    GTX1_RXUSRCLK2_IN                       : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX1_RXCDRRESET_IN                      : in   std_logic;
    GTX1_RXELECIDLE_OUT                     : out  std_logic;
    GTX1_RXEQMIX_IN                         : in   std_logic_vector(2 downto 0);
    GTX1_RXN_IN                             : in   std_logic;
    GTX1_RXP_IN                             : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GTX1_RXBUFRESET_IN                      : in   std_logic;
    GTX1_RXBUFSTATUS_OUT                    : out  std_logic_vector(2 downto 0);
    GTX1_RXCHANISALIGNED_OUT                : out  std_logic;
    GTX1_RXCHANREALIGN_OUT                  : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    GTX1_RXLOSSOFSYNC_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTX1_GTXRXRESET_IN                      : in   std_logic;
    GTX1_MGTREFCLKRX_IN                     : in   std_logic;
    GTX1_PLLRXRESET_IN                      : in   std_logic;
    GTX1_RXPLLLKDET_OUT                     : out  std_logic;
    GTX1_RXRESETDONE_OUT                    : out  std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    GTX1_DADDR_IN                           : in   std_logic_vector(7 downto 0);
    GTX1_DCLK_IN                            : in   std_logic;
    GTX1_DEN_IN                             : in   std_logic;
    GTX1_DI_IN                              : in   std_logic_vector(15 downto 0);
    GTX1_DRDY_OUT                           : out  std_logic;
    GTX1_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GTX1_DWE_IN                             : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX1_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX1_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    GTX1_TXOUTCLK_OUT                       : out  std_logic;
    GTX1_TXRESET_IN                         : in   std_logic;
    GTX1_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX1_TXDIFFCTRL_IN                      : in   std_logic_vector(3 downto 0);
    GTX1_TXN_OUT                            : out  std_logic;
    GTX1_TXP_OUT                            : out  std_logic;
    GTX1_TXPOSTEMPHASIS_IN                  : in   std_logic_vector(4 downto 0);
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    GTX1_TXPREEMPHASIS_IN                   : in   std_logic_vector(3 downto 0);
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    GTX1_TXDLYALIGNDISABLE_IN               : in   std_logic;
    GTX1_TXDLYALIGNMONENB_IN                : in   std_logic;
    GTX1_TXDLYALIGNMONITOR_OUT              : out  std_logic_vector(7 downto 0);
    GTX1_TXDLYALIGNRESET_IN                 : in   std_logic;
    GTX1_TXENPMAPHASEALIGN_IN               : in   std_logic;
    GTX1_TXPMASETPHASE_IN                   : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX1_GTXTXRESET_IN                      : in   std_logic;
    GTX1_TXRESETDONE_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GTX1_TXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX1_TXPRBSFORCEERR_IN                  : in   std_logic;    
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GTX1_TXELECIDLE_IN                      : in   std_logic;



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX2  (X0Y2)

    ------------------------ Loopback and Powerdown Ports ----------------------
    GTX2_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    GTX2_RXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    GTX2_TXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GTX2_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GTX2_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    GTX2_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GTX2_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GTX2_RXCHANBONDSEQ_OUT                  : out  std_logic;
    GTX2_RXCHBONDI_IN                       : in   std_logic_vector(3 downto 0);
    GTX2_RXCHBONDLEVEL_IN                   : in   std_logic_vector(2 downto 0);
    GTX2_RXCHBONDMASTER_IN                  : in   std_logic;
    GTX2_RXCHBONDO_OUT                      : out  std_logic_vector(3 downto 0);
    GTX2_RXCHBONDSLAVE_IN                   : in   std_logic;
    GTX2_RXENCHANSYNC_IN                    : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GTX2_RXCLKCORCNT_OUT                    : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GTX2_RXBYTEISALIGNED_OUT                : out  std_logic;
    GTX2_RXBYTEREALIGN_OUT                  : out  std_logic;
    GTX2_RXCOMMADET_OUT                     : out  std_logic;
    GTX2_RXENMCOMMAALIGN_IN                 : in   std_logic;
    GTX2_RXENPCOMMAALIGN_IN                 : in   std_logic;
    ----------------------- Receive Ports - PRBS Detection ---------------------
    GTX2_PRBSCNTRESET_IN                    : in   std_logic;
    GTX2_RXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX2_RXPRBSERR_OUT                      : out  std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTX2_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    GTX2_RXRESET_IN                         : in   std_logic;
    GTX2_RXUSRCLK2_IN                       : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX2_RXCDRRESET_IN                      : in   std_logic;
    GTX2_RXELECIDLE_OUT                     : out  std_logic;
    GTX2_RXEQMIX_IN                         : in   std_logic_vector(2 downto 0);
    GTX2_RXN_IN                             : in   std_logic;
    GTX2_RXP_IN                             : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GTX2_RXBUFRESET_IN                      : in   std_logic;
    GTX2_RXBUFSTATUS_OUT                    : out  std_logic_vector(2 downto 0);
    GTX2_RXCHANISALIGNED_OUT                : out  std_logic;
    GTX2_RXCHANREALIGN_OUT                  : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    GTX2_RXLOSSOFSYNC_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTX2_GTXRXRESET_IN                      : in   std_logic;
    GTX2_MGTREFCLKRX_IN                     : in   std_logic;
    GTX2_PLLRXRESET_IN                      : in   std_logic;
    GTX2_RXPLLLKDET_OUT                     : out  std_logic;
    GTX2_RXRESETDONE_OUT                    : out  std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    GTX2_DADDR_IN                           : in   std_logic_vector(7 downto 0);
    GTX2_DCLK_IN                            : in   std_logic;
    GTX2_DEN_IN                             : in   std_logic;
    GTX2_DI_IN                              : in   std_logic_vector(15 downto 0);
    GTX2_DRDY_OUT                           : out  std_logic;
    GTX2_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GTX2_DWE_IN                             : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX2_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX2_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    GTX2_TXOUTCLK_OUT                       : out  std_logic;
    GTX2_TXRESET_IN                         : in   std_logic;
    GTX2_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX2_TXDIFFCTRL_IN                      : in   std_logic_vector(3 downto 0);
    GTX2_TXN_OUT                            : out  std_logic;
    GTX2_TXP_OUT                            : out  std_logic;
    GTX2_TXPOSTEMPHASIS_IN                  : in   std_logic_vector(4 downto 0);
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    GTX2_TXPREEMPHASIS_IN                   : in   std_logic_vector(3 downto 0);
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    GTX2_TXDLYALIGNDISABLE_IN               : in   std_logic;
    GTX2_TXDLYALIGNMONENB_IN                : in   std_logic;
    GTX2_TXDLYALIGNMONITOR_OUT              : out  std_logic_vector(7 downto 0);
    GTX2_TXDLYALIGNRESET_IN                 : in   std_logic;
    GTX2_TXENPMAPHASEALIGN_IN               : in   std_logic;
    GTX2_TXPMASETPHASE_IN                   : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX2_GTXTXRESET_IN                      : in   std_logic;
    GTX2_TXRESETDONE_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GTX2_TXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX2_TXPRBSFORCEERR_IN                  : in   std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GTX2_TXELECIDLE_IN                      : in   std_logic;


    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX3  (X0Y3)

    ------------------------ Loopback and Powerdown Ports ----------------------
    GTX3_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    GTX3_RXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    GTX3_TXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GTX3_RXCHARISCOMMA_OUT                  : out  std_logic_vector(1 downto 0);
    GTX3_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    GTX3_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GTX3_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GTX3_RXCHANBONDSEQ_OUT                  : out  std_logic;
    GTX3_RXCHBONDI_IN                       : in   std_logic_vector(3 downto 0);
    GTX3_RXCHBONDLEVEL_IN                   : in   std_logic_vector(2 downto 0);
    GTX3_RXCHBONDMASTER_IN                  : in   std_logic;
    GTX3_RXCHBONDO_OUT                      : out  std_logic_vector(3 downto 0);
    GTX3_RXCHBONDSLAVE_IN                   : in   std_logic;
    GTX3_RXENCHANSYNC_IN                    : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GTX3_RXCLKCORCNT_OUT                    : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GTX3_RXBYTEISALIGNED_OUT                : out  std_logic;
    GTX3_RXBYTEREALIGN_OUT                  : out  std_logic;
    GTX3_RXCOMMADET_OUT                     : out  std_logic;
    GTX3_RXENMCOMMAALIGN_IN                 : in   std_logic;
    GTX3_RXENPCOMMAALIGN_IN                 : in   std_logic;
     ----------------------- Receive Ports - PRBS Detection ---------------------
    GTX3_PRBSCNTRESET_IN                    : in   std_logic;
    GTX3_RXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX3_RXPRBSERR_OUT                      : out  std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTX3_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    GTX3_RXRESET_IN                         : in   std_logic;
    GTX3_RXUSRCLK2_IN                       : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX3_RXCDRRESET_IN                      : in   std_logic;
    GTX3_RXELECIDLE_OUT                     : out  std_logic;
    GTX3_RXEQMIX_IN                         : in   std_logic_vector(2 downto 0);
    GTX3_RXN_IN                             : in   std_logic;
    GTX3_RXP_IN                             : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GTX3_RXBUFRESET_IN                      : in   std_logic;
    GTX3_RXBUFSTATUS_OUT                    : out  std_logic_vector(2 downto 0);
    GTX3_RXCHANISALIGNED_OUT                : out  std_logic;
    GTX3_RXCHANREALIGN_OUT                  : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    GTX3_RXLOSSOFSYNC_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTX3_GTXRXRESET_IN                      : in   std_logic;
    GTX3_MGTREFCLKRX_IN                     : in   std_logic;
    GTX3_PLLRXRESET_IN                      : in   std_logic;
    GTX3_RXPLLLKDET_OUT                     : out  std_logic;
    GTX3_RXRESETDONE_OUT                    : out  std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    GTX3_DADDR_IN                           : in   std_logic_vector(7 downto 0);
    GTX3_DCLK_IN                            : in   std_logic;
    GTX3_DEN_IN                             : in   std_logic;
    GTX3_DI_IN                              : in   std_logic_vector(15 downto 0);
    GTX3_DRDY_OUT                           : out  std_logic;
    GTX3_DRPDO_OUT                          : out  std_logic_vector(15 downto 0);
    GTX3_DWE_IN                             : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX3_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX3_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    GTX3_TXOUTCLK_OUT                       : out  std_logic;
    GTX3_TXRESET_IN                         : in   std_logic;
    GTX3_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX3_TXDIFFCTRL_IN                      : in   std_logic_vector(3 downto 0);
    GTX3_TXN_OUT                            : out  std_logic;
    GTX3_TXP_OUT                            : out  std_logic;
    GTX3_TXPOSTEMPHASIS_IN                  : in   std_logic_vector(4 downto 0);
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    GTX3_TXPREEMPHASIS_IN                   : in   std_logic_vector(3 downto 0);
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    GTX3_TXDLYALIGNDISABLE_IN               : in   std_logic;
    GTX3_TXDLYALIGNMONENB_IN                : in   std_logic;
    GTX3_TXDLYALIGNMONITOR_OUT              : out  std_logic_vector(7 downto 0);
    GTX3_TXDLYALIGNRESET_IN                 : in   std_logic;
    GTX3_TXENPMAPHASEALIGN_IN               : in   std_logic;
    GTX3_TXPMASETPHASE_IN                   : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX3_GTXTXRESET_IN                      : in   std_logic;
    GTX3_TXRESETDONE_OUT                    : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    GTX3_TXENPRBSTST_IN                     : in   std_logic_vector(2 downto 0);
    GTX3_TXPRBSFORCEERR_IN                  : in   std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GTX3_TXELECIDLE_IN                      : in   std_logic



);

    

end GTX_WRAPPER;

architecture RTL of GTX_WRAPPER is

attribute CORE_GENERATION_INFO : string;
attribute CORE_GENERATION_INFO of RTL : architecture is "GTX_WRAPPER,v6_gtxwizard_v1_5,{protocol_file=xaui}";
--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;

    signal  gtx0_share_rxpll_i           :   std_logic_vector(1 downto 0);
    signal  gtx0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);

    signal  gtx1_share_rxpll_i           :   std_logic_vector(1 downto 0);
    signal  gtx1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);

    signal  gtx2_share_rxpll_i           :   std_logic_vector(1 downto 0);
    signal  gtx2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);

    signal  gtx3_share_rxpll_i           :   std_logic_vector(1 downto 0);
    signal  gtx3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);

--*************************** Component Declarations **************************
component GTX_WRAPPER_GTX
generic
(
    -- Simulation attributes
    GTX_SIM_GTXRESET_SPEEDUP    : integer    := 0;

    -- Share RX PLL parameter
    GTX_TX_CLK_SOURCE           : string     := "TXPLL";
    -- Save power parameter
    GTX_POWER_SAVE              : bit_vector := "0000000000"
);
port
(
    ------------------------ Loopback and Powerdown Ports ----------------------
    LOOPBACK_IN                             : in   std_logic_vector(2 downto 0);
    RXPOWERDOWN_IN                          : in   std_logic_vector(1 downto 0);
    TXPOWERDOWN_IN                          : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISCOMMA_OUT                       : out  std_logic_vector(1 downto 0);
    RXCHARISK_OUT                           : out  std_logic_vector(1 downto 0);
    RXDISPERR_OUT                           : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    RXCHANBONDSEQ_OUT                       : out  std_logic;
    RXCHBONDI_IN                            : in   std_logic_vector(3 downto 0);
    RXCHBONDLEVEL_IN                        : in   std_logic_vector(2 downto 0);
    RXCHBONDMASTER_IN                       : in   std_logic;
    RXCHBONDO_OUT                           : out  std_logic_vector(3 downto 0);
    RXCHBONDSLAVE_IN                        : in   std_logic;
    RXENCHANSYNC_IN                         : in   std_logic;
     ------------------- Receive Ports - Clock Correction Ports -----------------
    RXCLKCORCNT_OUT                         : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXBYTEISALIGNED_OUT                     : out  std_logic;
    RXBYTEREALIGN_OUT                       : out  std_logic;
    RXCOMMADET_OUT                          : out  std_logic;
    RXENMCOMMAALIGN_IN                      : in   std_logic;
    RXENPCOMMAALIGN_IN                      : in   std_logic;
   ----------------------- Receive Ports - PRBS Detection ---------------------
    PRBSCNTRESET_IN                         : in   std_logic;
    RXENPRBSTST_IN                          : in   std_logic_vector(2 downto 0);
    RXPRBSERR_OUT                           : out  std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    RXDATA_OUT                              : out  std_logic_vector(15 downto 0);
    RXRESET_IN                              : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    RXCDRRESET_IN                           : in   std_logic;
    RXELECIDLE_OUT                          : out  std_logic;
    RXEQMIX_IN                              : in   std_logic_vector(2 downto 0);
    RXN_IN                                  : in   std_logic;
    RXP_IN                                  : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    RXBUFRESET_IN                           : in   std_logic;
    RXBUFSTATUS_OUT                         : out  std_logic_vector(2 downto 0);
    RXCHANISALIGNED_OUT                     : out  std_logic;
    RXCHANREALIGN_OUT                       : out  std_logic;
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    RXLOSSOFSYNC_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTXRXRESET_IN                           : in   std_logic;
    MGTREFCLKRX_IN                          : in   std_logic_vector(1 downto 0);
    PLLRXRESET_IN                           : in   std_logic;
    RXPLLLKDET_OUT                          : out  std_logic;
    RXRESETDONE_OUT                         : out  std_logic;
    ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
    DADDR_IN                                : in   std_logic_vector(7 downto 0);
    DCLK_IN                                 : in   std_logic;
    DEN_IN                                  : in   std_logic;
    DI_IN                                   : in   std_logic_vector(15 downto 0);
    DRDY_OUT                                : out  std_logic;
    DRPDO_OUT                               : out  std_logic_vector(15 downto 0);
    DWE_IN                                  : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TXCHARISK_IN                            : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA_IN                               : in   std_logic_vector(15 downto 0);
    TXOUTCLK_OUT                            : out  std_logic;
    TXRESET_IN                              : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    TXDIFFCTRL_IN                           : in   std_logic_vector(3 downto 0);
    TXN_OUT                                 : out  std_logic;
    TXP_OUT                                 : out  std_logic;
    TXPOSTEMPHASIS_IN                       : in   std_logic_vector(4 downto 0);
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TXPREEMPHASIS_IN                        : in   std_logic_vector(3 downto 0);
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    TXDLYALIGNDISABLE_IN                    : in   std_logic;
    TXDLYALIGNMONENB_IN                     : in   std_logic;
    TXDLYALIGNMONITOR_OUT                   : out  std_logic_vector(7 downto 0);
    TXDLYALIGNRESET_IN                      : in   std_logic;
    TXENPMAPHASEALIGN_IN                    : in   std_logic;
    TXPMASETPHASE_IN                        : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTXTXRESET_IN                           : in   std_logic;
    MGTREFCLKTX_IN                          : in   std_logic_vector(1 downto 0);
    PLLTXRESET_IN                           : in   std_logic;
    TXPLLLKDET_OUT                          : out  std_logic;
    TXRESETDONE_OUT                         : out  std_logic;
    --------------------- Transmit Ports - TX PRBS Generator -------------------
    TXENPRBSTST_IN                          : in   std_logic_vector(2 downto 0);
    TXPRBSFORCEERR_IN                       : in   std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TXELECIDLE_IN                           : in   std_logic



);
end component;

--********************************* Main Body of Code**************************

begin

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';

    gtx0_mgtrefclkrx_i <= (tied_to_ground_i & GTX0_MGTREFCLKRX_IN);
    gtx1_mgtrefclkrx_i <= (tied_to_ground_i & GTX1_MGTREFCLKRX_IN);
    gtx2_mgtrefclkrx_i <= (tied_to_ground_i & GTX2_MGTREFCLKRX_IN);
    gtx3_mgtrefclkrx_i <= (tied_to_ground_i & GTX3_MGTREFCLKRX_IN);


    --------------------------- GTX Instances  -------------------------------


    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX0  (X0Y0)

    gtx0_gtx_wrapper_i : GTX_WRAPPER_GTX
    generic map
    (
        -- Simulation attributes
        GTX_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,

        -- Share RX PLL parameter
        GTX_TX_CLK_SOURCE           => "RXPLL",
        -- Save power parameter
        GTX_POWER_SAVE              => "0000110100"
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GTX0_LOOPBACK_IN,
        RXPOWERDOWN_IN                  =>      GTX0_RXPOWERDOWN_IN,
        TXPOWERDOWN_IN                  =>      GTX0_TXPOWERDOWN_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GTX0_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GTX0_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GTX0_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GTX0_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GTX0_RXCHANBONDSEQ_OUT,
        RXCHBONDI_IN                    =>      GTX0_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GTX0_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GTX0_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GTX0_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GTX0_RXCHBONDSLAVE_IN,
        RXENCHANSYNC_IN                 =>      GTX0_RXENCHANSYNC_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GTX0_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GTX0_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GTX0_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GTX0_RXCOMMADET_OUT,
        RXENMCOMMAALIGN_IN              =>      GTX0_RXENMCOMMAALIGN_IN,
        RXENPCOMMAALIGN_IN              =>      GTX0_RXENPCOMMAALIGN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        PRBSCNTRESET_IN                 =>      GTX0_PRBSCNTRESET_IN,
        RXENPRBSTST_IN                  =>      GTX0_RXENPRBSTST_IN,
        RXPRBSERR_OUT                   =>      GTX0_RXPRBSERR_OUT,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA_OUT                      =>      GTX0_RXDATA_OUT,
        RXRESET_IN                      =>      GTX0_RXRESET_IN,
        RXUSRCLK2_IN                    =>      GTX0_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET_IN                   =>      GTX0_RXCDRRESET_IN,
        RXELECIDLE_OUT                  =>      GTX0_RXELECIDLE_OUT,
        RXEQMIX_IN                      =>      GTX0_RXEQMIX_IN,
        RXN_IN                          =>      GTX0_RXN_IN,
        RXP_IN                          =>      GTX0_RXP_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GTX0_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GTX0_RXBUFSTATUS_OUT,
        RXCHANISALIGNED_OUT             =>      GTX0_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GTX0_RXCHANREALIGN_OUT,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC_OUT                =>      GTX0_RXLOSSOFSYNC_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GTXRXRESET_IN                   =>      GTX0_GTXRXRESET_IN,
        MGTREFCLKRX_IN                  =>      gtx0_mgtrefclkrx_i,
        PLLRXRESET_IN                   =>      GTX0_PLLRXRESET_IN,
        RXPLLLKDET_OUT                  =>      GTX0_RXPLLLKDET_OUT,
        RXRESETDONE_OUT                 =>      GTX0_RXRESETDONE_OUT,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      GTX0_DADDR_IN,
        DCLK_IN                         =>      GTX0_DCLK_IN,
        DEN_IN                          =>      GTX0_DEN_IN,
        DI_IN                           =>      GTX0_DI_IN,
        DRDY_OUT                        =>      GTX0_DRDY_OUT,
        DRPDO_OUT                       =>      GTX0_DRPDO_OUT,
        DWE_IN                          =>      GTX0_DWE_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GTX0_TXCHARISK_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GTX0_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GTX0_TXOUTCLK_OUT,
        TXRESET_IN                      =>      GTX0_TXRESET_IN,
        TXUSRCLK2_IN                    =>      GTX0_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        TXDIFFCTRL_IN                   =>      GTX0_TXDIFFCTRL_IN,
        TXN_OUT                         =>      GTX0_TXN_OUT,
        TXP_OUT                         =>      GTX0_TXP_OUT,
        TXPOSTEMPHASIS_IN               =>      GTX0_TXPOSTEMPHASIS_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXPREEMPHASIS_IN                =>      GTX0_TXPREEMPHASIS_IN,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXDLYALIGNDISABLE_IN            =>      GTX0_TXDLYALIGNDISABLE_IN,
        TXDLYALIGNMONENB_IN             =>      GTX0_TXDLYALIGNMONENB_IN,
        TXDLYALIGNMONITOR_OUT           =>      GTX0_TXDLYALIGNMONITOR_OUT,
        TXDLYALIGNRESET_IN              =>      GTX0_TXDLYALIGNRESET_IN,
        TXENPMAPHASEALIGN_IN            =>      GTX0_TXENPMAPHASEALIGN_IN,
        TXPMASETPHASE_IN                =>      GTX0_TXPMASETPHASE_IN,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTXTXRESET_IN                   =>      GTX0_GTXTXRESET_IN,
        MGTREFCLKTX_IN                  =>      gtx0_mgtrefclkrx_i,
        PLLTXRESET_IN                   =>      tied_to_ground_i,
        TXPLLLKDET_OUT                  =>      open,
        TXRESETDONE_OUT                 =>      GTX0_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXENPRBSTST_IN                  =>      GTX0_TXENPRBSTST_IN,
        TXPRBSFORCEERR_IN               =>      GTX0_TXPRBSFORCEERR_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GTX0_TXELECIDLE_IN


    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX1  (X0Y1)

    gtx1_gtx_wrapper_i : GTX_WRAPPER_GTX
    generic map
    (
        -- Simulation attributes
        GTX_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,

        -- Share RX PLL parameter
        GTX_TX_CLK_SOURCE           => "RXPLL",
        -- Save power parameter
        GTX_POWER_SAVE              => "0000110100"
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GTX1_LOOPBACK_IN,
        RXPOWERDOWN_IN                  =>      GTX1_RXPOWERDOWN_IN,
        TXPOWERDOWN_IN                  =>      GTX1_TXPOWERDOWN_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GTX1_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GTX1_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GTX1_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GTX1_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GTX1_RXCHANBONDSEQ_OUT,
        RXCHBONDI_IN                    =>      GTX1_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GTX1_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GTX1_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GTX1_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GTX1_RXCHBONDSLAVE_IN,
        RXENCHANSYNC_IN                 =>      GTX1_RXENCHANSYNC_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GTX1_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GTX1_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GTX1_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GTX1_RXCOMMADET_OUT,
        RXENMCOMMAALIGN_IN              =>      GTX1_RXENMCOMMAALIGN_IN,
        RXENPCOMMAALIGN_IN              =>      GTX1_RXENPCOMMAALIGN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        PRBSCNTRESET_IN                 =>      GTX1_PRBSCNTRESET_IN,
        RXENPRBSTST_IN                  =>      GTX1_RXENPRBSTST_IN,
        RXPRBSERR_OUT                   =>      GTX1_RXPRBSERR_OUT,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA_OUT                      =>      GTX1_RXDATA_OUT,
        RXRESET_IN                      =>      GTX1_RXRESET_IN,
        RXUSRCLK2_IN                    =>      GTX1_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET_IN                   =>      GTX1_RXCDRRESET_IN,
        RXELECIDLE_OUT                  =>      GTX1_RXELECIDLE_OUT,
        RXEQMIX_IN                      =>      GTX1_RXEQMIX_IN,
        RXN_IN                          =>      GTX1_RXN_IN,
        RXP_IN                          =>      GTX1_RXP_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GTX1_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GTX1_RXBUFSTATUS_OUT,
        RXCHANISALIGNED_OUT             =>      GTX1_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GTX1_RXCHANREALIGN_OUT,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC_OUT                =>      GTX1_RXLOSSOFSYNC_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GTXRXRESET_IN                   =>      GTX1_GTXRXRESET_IN,
        MGTREFCLKRX_IN                  =>      gtx1_mgtrefclkrx_i,
        PLLRXRESET_IN                   =>      GTX1_PLLRXRESET_IN,
        RXPLLLKDET_OUT                  =>      GTX1_RXPLLLKDET_OUT,
        RXRESETDONE_OUT                 =>      GTX1_RXRESETDONE_OUT,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      GTX1_DADDR_IN,
        DCLK_IN                         =>      GTX1_DCLK_IN,
        DEN_IN                          =>      GTX1_DEN_IN,
        DI_IN                           =>      GTX1_DI_IN,
        DRDY_OUT                        =>      GTX1_DRDY_OUT,
        DRPDO_OUT                       =>      GTX1_DRPDO_OUT,
        DWE_IN                          =>      GTX1_DWE_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GTX1_TXCHARISK_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GTX1_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GTX1_TXOUTCLK_OUT,
        TXRESET_IN                      =>      GTX1_TXRESET_IN,
        TXUSRCLK2_IN                    =>      GTX1_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        TXDIFFCTRL_IN                   =>      GTX1_TXDIFFCTRL_IN,
        TXN_OUT                         =>      GTX1_TXN_OUT,
        TXP_OUT                         =>      GTX1_TXP_OUT,
        TXPOSTEMPHASIS_IN               =>      GTX1_TXPOSTEMPHASIS_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXPREEMPHASIS_IN                =>      GTX1_TXPREEMPHASIS_IN,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXDLYALIGNDISABLE_IN            =>      GTX1_TXDLYALIGNDISABLE_IN,
        TXDLYALIGNMONENB_IN             =>      GTX1_TXDLYALIGNMONENB_IN,
        TXDLYALIGNMONITOR_OUT           =>      GTX1_TXDLYALIGNMONITOR_OUT,
        TXDLYALIGNRESET_IN              =>      GTX1_TXDLYALIGNRESET_IN,
        TXENPMAPHASEALIGN_IN            =>      GTX1_TXENPMAPHASEALIGN_IN,
        TXPMASETPHASE_IN                =>      GTX1_TXPMASETPHASE_IN,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTXTXRESET_IN                   =>      GTX1_GTXTXRESET_IN,
        MGTREFCLKTX_IN                  =>      gtx1_mgtrefclkrx_i,
        PLLTXRESET_IN                   =>      tied_to_ground_i,
        TXPLLLKDET_OUT                  =>      open,
        TXRESETDONE_OUT                 =>      GTX1_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXENPRBSTST_IN                  =>      GTX1_TXENPRBSTST_IN,
        TXPRBSFORCEERR_IN               =>      GTX1_TXPRBSFORCEERR_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GTX1_TXELECIDLE_IN


    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX2  (X0Y2)

    gtx2_gtx_wrapper_i : GTX_WRAPPER_GTX
    generic map
    (
        -- Simulation attributes
        GTX_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,

        -- Share RX PLL parameter
        GTX_TX_CLK_SOURCE           => "RXPLL",
        -- Save power parameter
        GTX_POWER_SAVE              => "0000110100"
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GTX2_LOOPBACK_IN,
        RXPOWERDOWN_IN                  =>      GTX2_RXPOWERDOWN_IN,
        TXPOWERDOWN_IN                  =>      GTX2_TXPOWERDOWN_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GTX2_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GTX2_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GTX2_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GTX2_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GTX2_RXCHANBONDSEQ_OUT,
        RXCHBONDI_IN                    =>      GTX2_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GTX2_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GTX2_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GTX2_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GTX2_RXCHBONDSLAVE_IN,
        RXENCHANSYNC_IN                 =>      GTX2_RXENCHANSYNC_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GTX2_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GTX2_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GTX2_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GTX2_RXCOMMADET_OUT,
        RXENMCOMMAALIGN_IN              =>      GTX2_RXENMCOMMAALIGN_IN,
        RXENPCOMMAALIGN_IN              =>      GTX2_RXENPCOMMAALIGN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        PRBSCNTRESET_IN                 =>      GTX2_PRBSCNTRESET_IN,
        RXENPRBSTST_IN                  =>      GTX2_RXENPRBSTST_IN,
        RXPRBSERR_OUT                   =>      GTX2_RXPRBSERR_OUT,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA_OUT                      =>      GTX2_RXDATA_OUT,
        RXRESET_IN                      =>      GTX2_RXRESET_IN,
        RXUSRCLK2_IN                    =>      GTX2_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET_IN                   =>      GTX2_RXCDRRESET_IN,
        RXELECIDLE_OUT                  =>      GTX2_RXELECIDLE_OUT,
        RXEQMIX_IN                      =>      GTX2_RXEQMIX_IN,
        RXN_IN                          =>      GTX2_RXN_IN,
        RXP_IN                          =>      GTX2_RXP_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GTX2_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GTX2_RXBUFSTATUS_OUT,
        RXCHANISALIGNED_OUT             =>      GTX2_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GTX2_RXCHANREALIGN_OUT,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC_OUT                =>      GTX2_RXLOSSOFSYNC_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GTXRXRESET_IN                   =>      GTX2_GTXRXRESET_IN,
        MGTREFCLKRX_IN                  =>      gtx2_mgtrefclkrx_i,
        PLLRXRESET_IN                   =>      GTX2_PLLRXRESET_IN,
        RXPLLLKDET_OUT                  =>      GTX2_RXPLLLKDET_OUT,
        RXRESETDONE_OUT                 =>      GTX2_RXRESETDONE_OUT,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      GTX2_DADDR_IN,
        DCLK_IN                         =>      GTX2_DCLK_IN,
        DEN_IN                          =>      GTX2_DEN_IN,
        DI_IN                           =>      GTX2_DI_IN,
        DRDY_OUT                        =>      GTX2_DRDY_OUT,
        DRPDO_OUT                       =>      GTX2_DRPDO_OUT,
        DWE_IN                          =>      GTX2_DWE_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GTX2_TXCHARISK_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GTX2_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GTX2_TXOUTCLK_OUT,
        TXRESET_IN                      =>      GTX2_TXRESET_IN,
        TXUSRCLK2_IN                    =>      GTX2_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        TXDIFFCTRL_IN                   =>      GTX2_TXDIFFCTRL_IN,
        TXN_OUT                         =>      GTX2_TXN_OUT,
        TXP_OUT                         =>      GTX2_TXP_OUT,
        TXPOSTEMPHASIS_IN               =>      GTX2_TXPOSTEMPHASIS_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXPREEMPHASIS_IN                =>      GTX2_TXPREEMPHASIS_IN,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXDLYALIGNDISABLE_IN            =>      GTX2_TXDLYALIGNDISABLE_IN,
        TXDLYALIGNMONENB_IN             =>      GTX2_TXDLYALIGNMONENB_IN,
        TXDLYALIGNMONITOR_OUT           =>      GTX2_TXDLYALIGNMONITOR_OUT,
        TXDLYALIGNRESET_IN              =>      GTX2_TXDLYALIGNRESET_IN,
        TXENPMAPHASEALIGN_IN            =>      GTX2_TXENPMAPHASEALIGN_IN,
        TXPMASETPHASE_IN                =>      GTX2_TXPMASETPHASE_IN,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTXTXRESET_IN                   =>      GTX2_GTXTXRESET_IN,
        MGTREFCLKTX_IN                  =>      gtx2_mgtrefclkrx_i,
        PLLTXRESET_IN                   =>      tied_to_ground_i,
        TXPLLLKDET_OUT                  =>      open,
        TXRESETDONE_OUT                 =>      GTX2_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXENPRBSTST_IN                  =>      GTX2_TXENPRBSTST_IN,
        TXPRBSFORCEERR_IN               =>      GTX2_TXPRBSFORCEERR_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GTX2_TXELECIDLE_IN


    );



    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX3  (X0Y3)

    gtx3_gtx_wrapper_i : GTX_WRAPPER_GTX
    generic map
    (
        -- Simulation attributes
        GTX_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,

        -- Share RX PLL parameter
        GTX_TX_CLK_SOURCE           => "RXPLL",
        -- Save power parameter
        GTX_POWER_SAVE              => "0000110100"
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GTX3_LOOPBACK_IN,
        RXPOWERDOWN_IN                  =>      GTX3_RXPOWERDOWN_IN,
        TXPOWERDOWN_IN                  =>      GTX3_TXPOWERDOWN_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA_OUT               =>      GTX3_RXCHARISCOMMA_OUT,
        RXCHARISK_OUT                   =>      GTX3_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GTX3_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GTX3_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GTX3_RXCHANBONDSEQ_OUT,
        RXCHBONDI_IN                    =>      GTX3_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GTX3_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GTX3_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GTX3_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GTX3_RXCHBONDSLAVE_IN,
        RXENCHANSYNC_IN                 =>      GTX3_RXENCHANSYNC_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GTX3_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GTX3_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GTX3_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GTX3_RXCOMMADET_OUT,
        RXENMCOMMAALIGN_IN              =>      GTX3_RXENMCOMMAALIGN_IN,
        RXENPCOMMAALIGN_IN              =>      GTX3_RXENPCOMMAALIGN_IN,
        ----------------------- Receive Ports - PRBS Detection ---------------------
        PRBSCNTRESET_IN                 =>      GTX3_PRBSCNTRESET_IN,
        RXENPRBSTST_IN                  =>      GTX3_RXENPRBSTST_IN,
        RXPRBSERR_OUT                   =>      GTX3_RXPRBSERR_OUT,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA_OUT                      =>      GTX3_RXDATA_OUT,
        RXRESET_IN                      =>      GTX3_RXRESET_IN,
        RXUSRCLK2_IN                    =>      GTX3_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET_IN                   =>      GTX3_RXCDRRESET_IN,
        RXELECIDLE_OUT                  =>      GTX3_RXELECIDLE_OUT,
        RXEQMIX_IN                      =>      GTX3_RXEQMIX_IN,
        RXN_IN                          =>      GTX3_RXN_IN,
        RXP_IN                          =>      GTX3_RXP_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GTX3_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GTX3_RXBUFSTATUS_OUT,
        RXCHANISALIGNED_OUT             =>      GTX3_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GTX3_RXCHANREALIGN_OUT,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC_OUT                =>      GTX3_RXLOSSOFSYNC_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GTXRXRESET_IN                   =>      GTX3_GTXRXRESET_IN,
        MGTREFCLKRX_IN                  =>      gtx3_mgtrefclkrx_i,
        PLLRXRESET_IN                   =>      GTX3_PLLRXRESET_IN,
        RXPLLLKDET_OUT                  =>      GTX3_RXPLLLKDET_OUT,
        RXRESETDONE_OUT                 =>      GTX3_RXRESETDONE_OUT,
        ------------- Shared Ports - Dynamic Reconfiguration Port (DRP) ------------
        DADDR_IN                        =>      GTX3_DADDR_IN,
        DCLK_IN                         =>      GTX3_DCLK_IN,
        DEN_IN                          =>      GTX3_DEN_IN,
        DI_IN                           =>      GTX3_DI_IN,
        DRDY_OUT                        =>      GTX3_DRDY_OUT,
        DRPDO_OUT                       =>      GTX3_DRPDO_OUT,
        DWE_IN                          =>      GTX3_DWE_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARISK_IN                    =>      GTX3_TXCHARISK_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GTX3_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GTX3_TXOUTCLK_OUT,
        TXRESET_IN                      =>      GTX3_TXRESET_IN,
        TXUSRCLK2_IN                    =>      GTX3_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        TXDIFFCTRL_IN                   =>      GTX3_TXDIFFCTRL_IN,
        TXN_OUT                         =>      GTX3_TXN_OUT,
        TXP_OUT                         =>      GTX3_TXP_OUT,
        TXPOSTEMPHASIS_IN               =>      GTX3_TXPOSTEMPHASIS_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXPREEMPHASIS_IN                =>      GTX3_TXPREEMPHASIS_IN,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        TXDLYALIGNDISABLE_IN            =>      GTX3_TXDLYALIGNDISABLE_IN,
        TXDLYALIGNMONENB_IN             =>      GTX3_TXDLYALIGNMONENB_IN,
        TXDLYALIGNMONITOR_OUT           =>      GTX3_TXDLYALIGNMONITOR_OUT,
        TXDLYALIGNRESET_IN              =>      GTX3_TXDLYALIGNRESET_IN,
        TXENPMAPHASEALIGN_IN            =>      GTX3_TXENPMAPHASEALIGN_IN,
        TXPMASETPHASE_IN                =>      GTX3_TXPMASETPHASE_IN,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTXTXRESET_IN                   =>      GTX3_GTXTXRESET_IN,
        MGTREFCLKTX_IN                  =>      gtx3_mgtrefclkrx_i,
        PLLTXRESET_IN                   =>      tied_to_ground_i,
        TXPLLLKDET_OUT                  =>      open,
        TXRESETDONE_OUT                 =>      GTX3_TXRESETDONE_OUT,
        --------------------- Transmit Ports - TX PRBS Generator -------------------
        TXENPRBSTST_IN                  =>      GTX3_TXENPRBSTST_IN,
        TXPRBSFORCEERR_IN               =>      GTX3_TXPRBSFORCEERR_IN,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXELECIDLE_IN                   =>      GTX3_TXELECIDLE_IN

    );




end RTL;
