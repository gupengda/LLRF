-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.12
--  \   \         Application : Virtex-6 FPGA GTX Transceiver Wizard
--  /   /         Filename : v6_gtxwizard_v1_12.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module V6_GTXWIZARD_V1_12 (a GTX Wrapper)
-- Generated by Xilinx Virtex-6 FPGA GTX Transceiver Wizard
-- 
-- 
-- (c) Copyright 2009-2011 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity v6_gtxwizard_v1_12 is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset

    -- Reference Clock Frequency
    REF_CLK_FREQ                    : integer := 100
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX0  (X0Y0)
    
    ------------------------ Loopback and Powerdown Ports ----------------------
    GTX0_LOOPBACK_IN                        : in   std_logic_vector(2 downto 0);
    GTX0_RXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    GTX0_TXPOWERDOWN_IN                     : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    GTX0_RXCHARISK_OUT                      : out  std_logic_vector(1 downto 0);
    GTX0_RXDISPERR_OUT                      : out  std_logic_vector(1 downto 0);
    GTX0_RXNOTINTABLE_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    GTX0_RXCHANBONDSEQ_OUT                  : out  std_logic;
    GTX0_RXCHBONDI_IN                       : in   std_logic_vector(3 downto 0);
    GTX0_RXCHBONDLEVEL_IN                   : in   std_logic_vector(2 downto 0);
    GTX0_RXCHBONDMASTER_IN                  : in   std_logic;
    GTX0_RXCHBONDO_OUT                      : out  std_logic_vector(3 downto 0);
    GTX0_RXCHBONDSLAVE_IN                   : in   std_logic;
    GTX0_RXENCHANSYNC_IN                    : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    GTX0_RXCLKCORCNT_OUT                    : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    GTX0_RXBYTEISALIGNED_OUT                : out  std_logic;
    GTX0_RXBYTEREALIGN_OUT                  : out  std_logic;
    GTX0_RXCOMMADET_OUT                     : out  std_logic;
    GTX0_RXENMCOMMAALIGN_IN                 : in   std_logic;
    GTX0_RXENPCOMMAALIGN_IN                 : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    GTX0_RXDATA_OUT                         : out  std_logic_vector(15 downto 0);
    GTX0_RXRESET_IN                         : in   std_logic;
    GTX0_RXUSRCLK2_IN                       : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX0_RXCDRRESET_IN                      : in   std_logic;
    GTX0_RXELECIDLE_OUT                     : out  std_logic;
    GTX0_RXN_IN                             : in   std_logic;
    GTX0_RXP_IN                             : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    GTX0_RXBUFRESET_IN                      : in   std_logic;
    GTX0_RXBUFSTATUS_OUT                    : out  std_logic_vector(2 downto 0);
    GTX0_RXCHANISALIGNED_OUT                : out  std_logic;
    GTX0_RXCHANREALIGN_OUT                  : out  std_logic;
    GTX0_RXSTATUS_OUT                       : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    GTX0_RXLOSSOFSYNC_OUT                   : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTX0_GTXRXRESET_IN                      : in   std_logic;
    GTX0_MGTREFCLKRX_IN                     : in   std_logic;
    GTX0_PLLRXRESET_IN                      : in   std_logic;
    GTX0_RXPLLLKDET_OUT                     : out  std_logic;
    GTX0_RXRATE_IN                          : in   std_logic_vector(1 downto 0);
    GTX0_RXRATEDONE_OUT                     : out  std_logic;
    GTX0_RXRESETDONE_OUT                    : out  std_logic;
    -------------- Receive Ports - RX Pipe Control for PCI Express -------------
    GTX0_PHYSTATUS_OUT                      : out  std_logic;
    GTX0_RXVALID_OUT                        : out  std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GTX0_RXPOLARITY_IN                      : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX0_TXCHARDISPMODE_IN                  : in   std_logic_vector(1 downto 0);
    GTX0_TXCHARISK_IN                       : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX0_TXDATA_IN                          : in   std_logic_vector(15 downto 0);
    GTX0_TXOUTCLK_OUT                       : out  std_logic;
    GTX0_TXRESET_IN                         : in   std_logic;
    GTX0_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX0_TXN_OUT                            : out  std_logic;
    GTX0_TXP_OUT                            : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX0_GTXTXRESET_IN                      : in   std_logic;
    GTX0_MGTREFCLKTX_IN                     : in   std_logic;
    GTX0_PLLTXRESET_IN                      : in   std_logic;
    GTX0_TXPLLLKDET_OUT                     : out  std_logic;
    GTX0_TXRATE_IN                          : in   std_logic_vector(1 downto 0);
    GTX0_TXRATEDONE_OUT                     : out  std_logic;
    GTX0_TXRESETDONE_OUT                    : out  std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    GTX0_TXDEEMPH_IN                        : in   std_logic;
    GTX0_TXDETECTRX_IN                      : in   std_logic;
    GTX0_TXELECIDLE_IN                      : in   std_logic;
    GTX0_TXMARGIN_IN                        : in   std_logic_vector(2 downto 0);
    GTX0_TXPDOWNASYNCH_IN                   : in   std_logic;
    GTX0_TXSWING_IN                         : in   std_logic

    
);


end v6_gtxwizard_v1_12;
    
architecture RTL of v6_gtxwizard_v1_12 is

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "v6_gtxwizard_v1_12,v6_gtxwizard_v1_12,{protocol_file=pcie_gen2}";

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;


  
    signal  gtx0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
    signal  gtx0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
   
--*************************** Component Declarations **************************
component v6_gtxwizard_v1_12_gtx
generic
(
    -- Simulation attributes
    GTX_SIM_GTXRESET_SPEEDUP    : integer    := 0;
    
    -- Share RX PLL parameter
    GTX_TX_CLK_SOURCE           : string     := "TXPLL";
    -- Save power parameter
    GTX_POWER_SAVE              : bit_vector := "0000000000";

    -- Reference Clock Frequency
    REF_CLK_FREQ                    : integer := 100
);
port 
(   
    ------------------------ Loopback and Powerdown Ports ----------------------
    LOOPBACK_IN                             : in   std_logic_vector(2 downto 0);
    RXPOWERDOWN_IN                          : in   std_logic_vector(1 downto 0);
    TXPOWERDOWN_IN                          : in   std_logic_vector(1 downto 0);
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISK_OUT                           : out  std_logic_vector(1 downto 0);
    RXDISPERR_OUT                           : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------- Receive Ports - Channel Bonding Ports ------------------
    RXCHANBONDSEQ_OUT                       : out  std_logic;
    RXCHBONDI_IN                            : in   std_logic_vector(3 downto 0);
    RXCHBONDLEVEL_IN                        : in   std_logic_vector(2 downto 0);
    RXCHBONDMASTER_IN                       : in   std_logic;
    RXCHBONDO_OUT                           : out  std_logic_vector(3 downto 0);
    RXCHBONDSLAVE_IN                        : in   std_logic;
    RXENCHANSYNC_IN                         : in   std_logic;
    ------------------- Receive Ports - Clock Correction Ports -----------------
    RXCLKCORCNT_OUT                         : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXBYTEISALIGNED_OUT                     : out  std_logic;
    RXBYTEREALIGN_OUT                       : out  std_logic;
    RXCOMMADET_OUT                          : out  std_logic;
    RXENMCOMMAALIGN_IN                      : in   std_logic;
    RXENPCOMMAALIGN_IN                      : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    RXDATA_OUT                              : out  std_logic_vector(15 downto 0);
    RXRESET_IN                              : in   std_logic;
    RXUSRCLK2_IN                            : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    RXCDRRESET_IN                           : in   std_logic;
    RXELECIDLE_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic;
    RXP_IN                                  : in   std_logic;
    -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    RXBUFRESET_IN                           : in   std_logic;
    RXBUFSTATUS_OUT                         : out  std_logic_vector(2 downto 0);
    RXCHANISALIGNED_OUT                     : out  std_logic;
    RXCHANREALIGN_OUT                       : out  std_logic;
    RXSTATUS_OUT                            : out  std_logic_vector(2 downto 0);
    --------------- Receive Ports - RX Loss-of-sync State Machine --------------
    RXLOSSOFSYNC_OUT                        : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX PLL Ports ----------------------
    GTXRXRESET_IN                           : in   std_logic;
    MGTREFCLKRX_IN                          : in   std_logic_vector(1 downto 0);
    PLLRXRESET_IN                           : in   std_logic;
    RXPLLLKDET_OUT                          : out  std_logic;
    RXRATE_IN                               : in   std_logic_vector(1 downto 0);
    RXRATEDONE_OUT                          : out  std_logic;
    RXRESETDONE_OUT                         : out  std_logic;
    -------------- Receive Ports - RX Pipe Control for PCI Express -------------
    PHYSTATUS_OUT                           : out  std_logic;
    RXVALID_OUT                             : out  std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    RXPOLARITY_IN                           : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TXCHARDISPMODE_IN                       : in   std_logic_vector(1 downto 0);
    TXCHARISK_IN                            : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA_IN                               : in   std_logic_vector(15 downto 0);
    TXOUTCLK_OUT                            : out  std_logic;
    TXRESET_IN                              : in   std_logic;
    TXUSRCLK2_IN                            : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    TXN_OUT                                 : out  std_logic;
    TXP_OUT                                 : out  std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTXTXRESET_IN                           : in   std_logic;
    MGTREFCLKTX_IN                          : in   std_logic_vector(1 downto 0);
    PLLTXRESET_IN                           : in   std_logic;
    TXPLLLKDET_OUT                          : out  std_logic;
    TXRATE_IN                               : in   std_logic_vector(1 downto 0);
    TXRATEDONE_OUT                          : out  std_logic;
    TXRESETDONE_OUT                         : out  std_logic;
    ----------------- Transmit Ports - TX Ports for PCI Express ----------------
    TXDEEMPH_IN                             : in   std_logic;
    TXDETECTRX_IN                           : in   std_logic;
    TXELECIDLE_IN                           : in   std_logic;
    TXMARGIN_IN                             : in   std_logic_vector(2 downto 0);
    TXPDOWNASYNCH_IN                        : in   std_logic;
    TXSWING_IN                              : in   std_logic


);
end component;


--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
                     

   
    gtx0_mgtrefclktx_i <= (tied_to_ground_i & GTX0_MGTREFCLKTX_IN);
    gtx0_mgtrefclkrx_i <= (tied_to_ground_i & GTX0_MGTREFCLKRX_IN);

 
    --------------------------- GTX Instances  -------------------------------   


    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX0  (X0Y0)

    gtx0_v6_gtxwizard_v1_12_i : v6_gtxwizard_v1_12_gtx
    generic map
    (
        -- Simulation attributes
        GTX_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        
        -- Share RX PLL parameter
        GTX_TX_CLK_SOURCE           => "TXPLL",
        -- Save power parameter
        GTX_POWER_SAVE              => "0000110000",

        -- Tx/Rx PLL dividers
        REF_CLK_FREQ                => REF_CLK_FREQ
    )
    port map
    (
        ------------------------ Loopback and Powerdown Ports ----------------------
        LOOPBACK_IN                     =>      GTX0_LOOPBACK_IN,
        RXPOWERDOWN_IN                  =>      GTX0_RXPOWERDOWN_IN,
        TXPOWERDOWN_IN                  =>      GTX0_TXPOWERDOWN_IN,
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISK_OUT                   =>      GTX0_RXCHARISK_OUT,
        RXDISPERR_OUT                   =>      GTX0_RXDISPERR_OUT,
        RXNOTINTABLE_OUT                =>      GTX0_RXNOTINTABLE_OUT,
        ------------------- Receive Ports - Channel Bonding Ports ------------------
        RXCHANBONDSEQ_OUT               =>      GTX0_RXCHANBONDSEQ_OUT,
        RXCHBONDI_IN                    =>      GTX0_RXCHBONDI_IN,
        RXCHBONDLEVEL_IN                =>      GTX0_RXCHBONDLEVEL_IN,
        RXCHBONDMASTER_IN               =>      GTX0_RXCHBONDMASTER_IN,
        RXCHBONDO_OUT                   =>      GTX0_RXCHBONDO_OUT,
        RXCHBONDSLAVE_IN                =>      GTX0_RXCHBONDSLAVE_IN,
        RXENCHANSYNC_IN                 =>      GTX0_RXENCHANSYNC_IN,
        ------------------- Receive Ports - Clock Correction Ports -----------------
        RXCLKCORCNT_OUT                 =>      GTX0_RXCLKCORCNT_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED_OUT             =>      GTX0_RXBYTEISALIGNED_OUT,
        RXBYTEREALIGN_OUT               =>      GTX0_RXBYTEREALIGN_OUT,
        RXCOMMADET_OUT                  =>      GTX0_RXCOMMADET_OUT,
        RXENMCOMMAALIGN_IN              =>      GTX0_RXENMCOMMAALIGN_IN,
        RXENPCOMMAALIGN_IN              =>      GTX0_RXENPCOMMAALIGN_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA_OUT                      =>      GTX0_RXDATA_OUT,
        RXRESET_IN                      =>      GTX0_RXRESET_IN,
        RXUSRCLK2_IN                    =>      GTX0_RXUSRCLK2_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXCDRRESET_IN                   =>      GTX0_RXCDRRESET_IN,
        RXELECIDLE_OUT                  =>      GTX0_RXELECIDLE_OUT,
        RXN_IN                          =>      GTX0_RXN_IN,
        RXP_IN                          =>      GTX0_RXP_IN,
        -------- Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
        RXBUFRESET_IN                   =>      GTX0_RXBUFRESET_IN,
        RXBUFSTATUS_OUT                 =>      GTX0_RXBUFSTATUS_OUT,
        RXCHANISALIGNED_OUT             =>      GTX0_RXCHANISALIGNED_OUT,
        RXCHANREALIGN_OUT               =>      GTX0_RXCHANREALIGN_OUT,
        RXSTATUS_OUT                    =>      GTX0_RXSTATUS_OUT,
        --------------- Receive Ports - RX Loss-of-sync State Machine --------------
        RXLOSSOFSYNC_OUT                =>      GTX0_RXLOSSOFSYNC_OUT,
        ------------------------ Receive Ports - RX PLL Ports ----------------------
        GTXRXRESET_IN                   =>      GTX0_GTXRXRESET_IN,
        MGTREFCLKRX_IN                  =>      gtx0_mgtrefclkrx_i,
        PLLRXRESET_IN                   =>      GTX0_PLLRXRESET_IN,
        RXPLLLKDET_OUT                  =>      GTX0_RXPLLLKDET_OUT,
        RXRATE_IN                       =>      GTX0_RXRATE_IN,
        RXRATEDONE_OUT                  =>      GTX0_RXRATEDONE_OUT,
        RXRESETDONE_OUT                 =>      GTX0_RXRESETDONE_OUT,
        -------------- Receive Ports - RX Pipe Control for PCI Express -------------
        PHYSTATUS_OUT                   =>      GTX0_PHYSTATUS_OUT,
        RXVALID_OUT                     =>      GTX0_RXVALID_OUT,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        RXPOLARITY_IN                   =>      GTX0_RXPOLARITY_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TXCHARDISPMODE_IN               =>      GTX0_TXCHARDISPMODE_IN,
        TXCHARISK_IN                    =>      GTX0_TXCHARISK_IN,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA_IN                       =>      GTX0_TXDATA_IN,
        TXOUTCLK_OUT                    =>      GTX0_TXOUTCLK_OUT,
        TXRESET_IN                      =>      GTX0_TXRESET_IN,
        TXUSRCLK2_IN                    =>      GTX0_TXUSRCLK2_IN,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        TXN_OUT                         =>      GTX0_TXN_OUT,
        TXP_OUT                         =>      GTX0_TXP_OUT,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTXTXRESET_IN                   =>      GTX0_GTXTXRESET_IN,
        MGTREFCLKTX_IN                  =>      gtx0_mgtrefclktx_i,
        PLLTXRESET_IN                   =>      GTX0_PLLTXRESET_IN,
        TXPLLLKDET_OUT                  =>      GTX0_TXPLLLKDET_OUT,
        TXRATE_IN                       =>      GTX0_TXRATE_IN,
        TXRATEDONE_OUT                  =>      GTX0_TXRATEDONE_OUT,
        TXRESETDONE_OUT                 =>      GTX0_TXRESETDONE_OUT,
        ----------------- Transmit Ports - TX Ports for PCI Express ----------------
        TXDEEMPH_IN                     =>      GTX0_TXDEEMPH_IN,
        TXDETECTRX_IN                   =>      GTX0_TXDETECTRX_IN,
        TXELECIDLE_IN                   =>      GTX0_TXELECIDLE_IN,
        TXMARGIN_IN                     =>      GTX0_TXMARGIN_IN,
        TXPDOWNASYNCH_IN                =>      GTX0_TXPDOWNASYNCH_IN,
        TXSWING_IN                      =>      GTX0_TXSWING_IN

    );

  
  
    

     
end RTL;
